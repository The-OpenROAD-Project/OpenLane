magic
tech sky130A
magscale 1 2
timestamp 1636140361
<< checkpaint >>
rect -1309 -1311 5698 22869
<< locali >>
rect 4337 11329 4371 11345
rect 3542 11295 4337 11329
rect 4337 11279 4371 11295
rect 2775 11059 2809 11075
rect 2775 11009 2809 11025
rect 2908 10935 2942 10951
rect 2908 10885 2942 10901
rect 3041 10811 3075 10827
rect 3041 10761 3075 10777
rect 3353 10622 3387 10638
rect 3353 10572 3387 10588
rect 4337 9915 4371 9931
rect 3064 9881 4337 9915
rect 4337 9865 4371 9881
rect 2760 9170 2794 9186
rect 2760 9120 2794 9136
rect 2875 9170 2909 9186
rect 2875 9120 2909 9136
rect 4337 8501 4371 8517
rect 3064 8467 4337 8501
rect 4337 8451 4371 8467
rect 2808 8231 2842 8247
rect 2808 8181 2842 8197
rect 2908 7983 2942 7999
rect 2908 7933 2942 7949
rect 3228 7350 3262 7832
rect 4227 7794 4261 7810
rect 4227 7744 4261 7760
rect 3043 7316 3262 7350
rect 4337 7087 4371 7103
rect 3542 7053 4337 7087
rect 4337 7037 4371 7053
rect 3353 6380 3387 6396
rect 3353 6330 3387 6346
rect 3041 6191 3075 6207
rect 3041 6141 3075 6157
rect 2908 6067 2942 6083
rect 2908 6017 2942 6033
rect 2775 5943 2809 5959
rect 2775 5893 2809 5909
rect 4337 5673 4371 5689
rect 3542 5639 4337 5673
rect 4337 5623 4371 5639
rect 2760 5004 2794 5020
rect 2760 4954 2794 4970
rect 4275 4966 4309 4982
rect 4275 4916 4309 4932
rect 4337 4259 4371 4275
rect 3442 4225 4337 4259
rect 4337 4209 4371 4225
rect 3253 3536 3287 3552
rect 3253 3486 3287 3502
rect 2908 3363 2942 3379
rect 2908 3313 2942 3329
rect 2808 3115 2842 3131
rect 2808 3065 2842 3081
rect 4337 2845 4371 2861
rect 3442 2811 4337 2845
rect 4337 2795 4371 2811
rect 3025 2541 3210 2575
rect 2760 2176 2794 2192
rect 3025 2176 3059 2541
rect 3276 2327 3310 2343
rect 3276 2277 3310 2293
rect 2892 2142 3059 2176
rect 3621 2154 3655 2170
rect 2760 2126 2794 2142
rect 3621 2104 3655 2120
rect 4337 1431 4371 1447
rect 3810 1397 4337 1431
rect 4337 1381 4371 1397
rect 4275 724 4309 740
rect 2760 686 2794 702
rect 4275 674 4309 690
rect 2760 636 2794 652
rect 4337 17 4371 33
rect 4337 -33 4371 -17
<< viali >>
rect 4337 11295 4371 11329
rect 2775 11025 2809 11059
rect 2908 10901 2942 10935
rect 3041 10777 3075 10811
rect 3353 10588 3387 10622
rect 4337 9881 4371 9915
rect 2760 9136 2794 9170
rect 2875 9136 2909 9170
rect 4337 8467 4371 8501
rect 2808 8197 2842 8231
rect 2908 7949 2942 7983
rect 4227 7760 4261 7794
rect 4337 7053 4371 7087
rect 3353 6346 3387 6380
rect 3041 6157 3075 6191
rect 2908 6033 2942 6067
rect 2775 5909 2809 5943
rect 4337 5639 4371 5673
rect 2760 4970 2794 5004
rect 4275 4932 4309 4966
rect 4337 4225 4371 4259
rect 3253 3502 3287 3536
rect 2908 3329 2942 3363
rect 2808 3081 2842 3115
rect 4337 2811 4371 2845
rect 3276 2293 3310 2327
rect 2760 2142 2794 2176
rect 3621 2120 3655 2154
rect 4337 1397 4371 1431
rect 2760 652 2794 686
rect 4275 690 4309 724
rect 4337 -17 4371 17
<< metal1 >>
rect 4322 11286 4328 11338
rect 4380 11286 4386 11338
rect 2006 11016 2012 11068
rect 2064 11056 2070 11068
rect 2763 11059 2821 11065
rect 2763 11056 2775 11059
rect 2064 11028 2775 11056
rect 2064 11016 2070 11028
rect 2763 11025 2775 11028
rect 2809 11025 2821 11059
rect 2763 11019 2821 11025
rect 2090 10892 2096 10944
rect 2148 10932 2154 10944
rect 2896 10935 2954 10941
rect 2896 10932 2908 10935
rect 2148 10904 2908 10932
rect 2148 10892 2154 10904
rect 2896 10901 2908 10904
rect 2942 10901 2954 10935
rect 2896 10895 2954 10901
rect 2342 10768 2348 10820
rect 2400 10808 2406 10820
rect 3029 10811 3087 10817
rect 3029 10808 3041 10811
rect 2400 10780 3041 10808
rect 2400 10768 2406 10780
rect 3029 10777 3041 10780
rect 3075 10777 3087 10811
rect 3029 10771 3087 10777
rect 3338 10579 3344 10631
rect 3396 10579 3402 10631
rect 4322 9872 4328 9924
rect 4380 9872 4386 9924
rect 2006 9127 2012 9179
rect 2064 9167 2070 9179
rect 2748 9170 2806 9176
rect 2748 9167 2760 9170
rect 2064 9139 2760 9167
rect 2064 9127 2070 9139
rect 2748 9136 2760 9139
rect 2794 9136 2806 9170
rect 2748 9130 2806 9136
rect 2860 9127 2866 9179
rect 2918 9127 2924 9179
rect 4322 8458 4328 8510
rect 4380 8458 4386 8510
rect 2174 8188 2180 8240
rect 2232 8228 2238 8240
rect 2796 8231 2854 8237
rect 2796 8228 2808 8231
rect 2232 8200 2808 8228
rect 2232 8188 2238 8200
rect 2796 8197 2808 8200
rect 2842 8197 2854 8231
rect 2796 8191 2854 8197
rect 2006 7940 2012 7992
rect 2064 7980 2070 7992
rect 2896 7983 2954 7989
rect 2896 7980 2908 7983
rect 2064 7952 2908 7980
rect 2064 7940 2070 7952
rect 2896 7949 2908 7952
rect 2942 7949 2954 7983
rect 2896 7943 2954 7949
rect 4212 7751 4218 7803
rect 4270 7751 4276 7803
rect 171 7027 177 7079
rect 229 7067 235 7079
rect 2006 7067 2012 7079
rect 229 7039 2012 7067
rect 229 7027 235 7039
rect 2006 7027 2012 7039
rect 2064 7027 2070 7079
rect 4322 7044 4328 7096
rect 4380 7044 4386 7096
rect 3338 6337 3344 6389
rect 3396 6337 3402 6389
rect 2090 6148 2096 6200
rect 2148 6188 2154 6200
rect 3029 6191 3087 6197
rect 3029 6188 3041 6191
rect 2148 6160 3041 6188
rect 2148 6148 2154 6160
rect 3029 6157 3041 6160
rect 3075 6157 3087 6191
rect 3029 6151 3087 6157
rect 1922 6024 1928 6076
rect 1980 6064 1986 6076
rect 2896 6067 2954 6073
rect 2896 6064 2908 6067
rect 1980 6036 2908 6064
rect 1980 6024 1986 6036
rect 2896 6033 2908 6036
rect 2942 6033 2954 6067
rect 2896 6027 2954 6033
rect 2258 5900 2264 5952
rect 2316 5940 2322 5952
rect 2763 5943 2821 5949
rect 2763 5940 2775 5943
rect 2316 5912 2775 5940
rect 2316 5900 2322 5912
rect 2763 5909 2775 5912
rect 2809 5909 2821 5943
rect 2763 5903 2821 5909
rect 4322 5630 4328 5682
rect 4380 5630 4386 5682
rect 2090 4961 2096 5013
rect 2148 5001 2154 5013
rect 2748 5004 2806 5010
rect 2748 5001 2760 5004
rect 2148 4973 2760 5001
rect 2148 4961 2154 4973
rect 2748 4970 2760 4973
rect 2794 4970 2806 5004
rect 2748 4964 2806 4970
rect 4260 4923 4266 4975
rect 4318 4923 4324 4975
rect 351 4216 357 4268
rect 409 4256 415 4268
rect 2426 4256 2432 4268
rect 409 4228 2432 4256
rect 409 4216 415 4228
rect 2426 4216 2432 4228
rect 2484 4216 2490 4268
rect 4322 4216 4328 4268
rect 4380 4216 4386 4268
rect 3238 3493 3244 3545
rect 3296 3493 3302 3545
rect 2510 3320 2516 3372
rect 2568 3360 2574 3372
rect 2896 3363 2954 3369
rect 2896 3360 2908 3363
rect 2568 3332 2908 3360
rect 2568 3320 2574 3332
rect 2896 3329 2908 3332
rect 2942 3329 2954 3363
rect 2896 3323 2954 3329
rect 2426 3072 2432 3124
rect 2484 3112 2490 3124
rect 2796 3115 2854 3121
rect 2796 3112 2808 3115
rect 2484 3084 2808 3112
rect 2484 3072 2490 3084
rect 2796 3081 2808 3084
rect 2842 3081 2854 3115
rect 2796 3075 2854 3081
rect 4322 2802 4328 2854
rect 4380 2802 4386 2854
rect 3261 2284 3267 2336
rect 3319 2284 3325 2336
rect 2426 2133 2432 2185
rect 2484 2173 2490 2185
rect 2748 2176 2806 2182
rect 2748 2173 2760 2176
rect 2484 2145 2760 2173
rect 2484 2133 2490 2145
rect 2748 2142 2760 2145
rect 2794 2142 2806 2176
rect 2748 2136 2806 2142
rect 3606 2111 3612 2163
rect 3664 2111 3670 2163
rect 4322 1388 4328 1440
rect 4380 1388 4386 1440
rect 2745 643 2751 695
rect 2803 643 2809 695
rect 4260 681 4266 733
rect 4318 681 4324 733
rect 4322 -26 4328 26
rect 4380 -26 4386 26
<< via1 >>
rect 4328 11329 4380 11338
rect 4328 11295 4337 11329
rect 4337 11295 4371 11329
rect 4371 11295 4380 11329
rect 4328 11286 4380 11295
rect 2012 11016 2064 11068
rect 2096 10892 2148 10944
rect 2348 10768 2400 10820
rect 3344 10622 3396 10631
rect 3344 10588 3353 10622
rect 3353 10588 3387 10622
rect 3387 10588 3396 10622
rect 3344 10579 3396 10588
rect 4328 9915 4380 9924
rect 4328 9881 4337 9915
rect 4337 9881 4371 9915
rect 4371 9881 4380 9915
rect 4328 9872 4380 9881
rect 2012 9127 2064 9179
rect 2866 9170 2918 9179
rect 2866 9136 2875 9170
rect 2875 9136 2909 9170
rect 2909 9136 2918 9170
rect 2866 9127 2918 9136
rect 4328 8501 4380 8510
rect 4328 8467 4337 8501
rect 4337 8467 4371 8501
rect 4371 8467 4380 8501
rect 4328 8458 4380 8467
rect 2180 8188 2232 8240
rect 2012 7940 2064 7992
rect 4218 7794 4270 7803
rect 4218 7760 4227 7794
rect 4227 7760 4261 7794
rect 4261 7760 4270 7794
rect 4218 7751 4270 7760
rect 177 7027 229 7079
rect 2012 7027 2064 7079
rect 4328 7087 4380 7096
rect 4328 7053 4337 7087
rect 4337 7053 4371 7087
rect 4371 7053 4380 7087
rect 4328 7044 4380 7053
rect 3344 6380 3396 6389
rect 3344 6346 3353 6380
rect 3353 6346 3387 6380
rect 3387 6346 3396 6380
rect 3344 6337 3396 6346
rect 2096 6148 2148 6200
rect 1928 6024 1980 6076
rect 2264 5900 2316 5952
rect 4328 5673 4380 5682
rect 4328 5639 4337 5673
rect 4337 5639 4371 5673
rect 4371 5639 4380 5673
rect 4328 5630 4380 5639
rect 2096 4961 2148 5013
rect 4266 4966 4318 4975
rect 4266 4932 4275 4966
rect 4275 4932 4309 4966
rect 4309 4932 4318 4966
rect 4266 4923 4318 4932
rect 357 4216 409 4268
rect 2432 4216 2484 4268
rect 4328 4259 4380 4268
rect 4328 4225 4337 4259
rect 4337 4225 4371 4259
rect 4371 4225 4380 4259
rect 4328 4216 4380 4225
rect 3244 3536 3296 3545
rect 3244 3502 3253 3536
rect 3253 3502 3287 3536
rect 3287 3502 3296 3536
rect 3244 3493 3296 3502
rect 2516 3320 2568 3372
rect 2432 3072 2484 3124
rect 4328 2845 4380 2854
rect 4328 2811 4337 2845
rect 4337 2811 4371 2845
rect 4371 2811 4380 2845
rect 4328 2802 4380 2811
rect 3267 2327 3319 2336
rect 3267 2293 3276 2327
rect 3276 2293 3310 2327
rect 3310 2293 3319 2327
rect 3267 2284 3319 2293
rect 2432 2133 2484 2185
rect 3612 2154 3664 2163
rect 3612 2120 3621 2154
rect 3621 2120 3655 2154
rect 3655 2120 3664 2154
rect 3612 2111 3664 2120
rect 4328 1431 4380 1440
rect 4328 1397 4337 1431
rect 4337 1397 4371 1431
rect 4371 1397 4380 1431
rect 4328 1388 4380 1397
rect 2751 686 2803 695
rect 2751 652 2760 686
rect 2760 652 2794 686
rect 2794 652 2803 686
rect 2751 643 2803 652
rect 4266 724 4318 733
rect 4266 690 4275 724
rect 4275 690 4309 724
rect 4309 690 4318 724
rect 4266 681 4318 690
rect 4328 17 4380 26
rect 4328 -17 4337 17
rect 4337 -17 4371 17
rect 4371 -17 4380 17
rect 4328 -26 4380 -17
<< metal2 >>
rect 1748 11472 1776 11994
rect 189 7085 217 11472
rect 1940 8624 1968 11388
rect 2024 11074 2052 11388
rect 2012 11068 2064 11074
rect 2012 11010 2064 11016
rect 2024 9185 2052 11010
rect 2108 10950 2136 11388
rect 2096 10944 2148 10950
rect 2096 10886 2148 10892
rect 2012 9179 2064 9185
rect 2012 9121 2064 9127
rect 1926 8615 1982 8624
rect 1926 8550 1982 8559
rect 177 7079 229 7085
rect 177 7021 229 7027
rect 1940 6082 1968 8550
rect 2024 7998 2052 9121
rect 2012 7992 2064 7998
rect 2012 7934 2064 7940
rect 2024 7085 2052 7934
rect 2012 7079 2064 7085
rect 2012 7021 2064 7027
rect 1928 6076 1980 6082
rect 1928 6018 1980 6024
rect 357 4268 409 4274
rect 357 4210 409 4216
rect 369 2828 397 4210
rect 1842 2351 1898 2360
rect 137 2238 203 2290
rect 1842 2286 1898 2295
rect 1498 1964 1554 1973
rect 1498 1899 1554 1908
rect 1498 920 1554 929
rect 1498 855 1554 864
rect 137 538 203 590
rect 1940 0 1968 6018
rect 2024 0 2052 7021
rect 2108 6206 2136 10886
rect 2192 8246 2220 11388
rect 2180 8240 2232 8246
rect 2180 8182 2232 8188
rect 2096 6200 2148 6206
rect 2096 6142 2148 6148
rect 2108 5019 2136 6142
rect 2096 5013 2148 5019
rect 2096 4955 2148 4961
rect 2108 1608 2136 4955
rect 2192 3556 2220 8182
rect 2276 5958 2304 11388
rect 2360 10826 2388 11388
rect 2348 10820 2400 10826
rect 2348 10762 2400 10768
rect 2264 5952 2316 5958
rect 2264 5894 2316 5900
rect 2178 3547 2234 3556
rect 2178 3482 2234 3491
rect 2094 1599 2150 1608
rect 2094 1534 2150 1543
rect 2108 0 2136 1534
rect 2192 0 2220 3482
rect 2276 1973 2304 5894
rect 2360 2360 2388 10762
rect 2444 4274 2472 11388
rect 2432 4268 2484 4274
rect 2432 4210 2484 4216
rect 2444 3130 2472 4210
rect 2528 3378 2556 11388
rect 4326 11340 4382 11349
rect 4326 11275 4382 11284
rect 3344 10631 3396 10637
rect 3396 10591 4438 10619
rect 3344 10573 3396 10579
rect 4326 9926 4382 9935
rect 4326 9861 4382 9870
rect 2866 9179 2918 9185
rect 2866 9121 2918 9127
rect 2878 8624 2906 9121
rect 2864 8615 2920 8624
rect 2864 8550 2920 8559
rect 4326 8512 4382 8521
rect 4326 8447 4382 8456
rect 4218 7803 4270 7809
rect 4270 7763 4438 7791
rect 4218 7745 4270 7751
rect 4326 7098 4382 7107
rect 4326 7033 4382 7042
rect 3344 6389 3396 6395
rect 3396 6349 4438 6377
rect 3344 6331 3396 6337
rect 4326 5684 4382 5693
rect 4326 5619 4382 5628
rect 4266 4975 4318 4981
rect 4318 4935 4438 4963
rect 4266 4917 4318 4923
rect 4326 4270 4382 4279
rect 4326 4205 4382 4214
rect 3242 3547 3298 3556
rect 3242 3482 3298 3491
rect 2516 3372 2568 3378
rect 2516 3314 2568 3320
rect 2432 3124 2484 3130
rect 2432 3066 2484 3072
rect 2346 2351 2402 2360
rect 2346 2286 2402 2295
rect 2262 1964 2318 1973
rect 2262 1899 2318 1908
rect 2276 0 2304 1899
rect 2360 0 2388 2286
rect 2444 2191 2472 3066
rect 2528 2347 2556 3314
rect 4326 2856 4382 2865
rect 4326 2791 4382 2800
rect 2514 2338 2570 2347
rect 2514 2273 2570 2282
rect 3265 2338 3321 2347
rect 3265 2273 3321 2282
rect 2432 2185 2484 2191
rect 2432 2127 2484 2133
rect 2444 178 2472 2127
rect 2528 929 2556 2273
rect 3612 2163 3664 2169
rect 3612 2105 3664 2111
rect 3624 1608 3652 2105
rect 3610 1599 3666 1608
rect 3610 1534 3666 1543
rect 4326 1442 4382 1451
rect 4326 1377 4382 1386
rect 2514 920 2570 929
rect 2514 855 2570 864
rect 2430 169 2486 178
rect 2430 104 2486 113
rect 2444 0 2472 104
rect 2528 0 2556 855
rect 4266 733 4318 739
rect 2751 695 2803 701
rect 4318 693 4438 721
rect 4266 675 4318 681
rect 2751 637 2803 643
rect 4278 178 4306 675
rect 4264 169 4320 178
rect 4264 104 4320 113
rect 4326 28 4382 37
rect 4326 -37 4382 -28
<< via2 >>
rect 1926 8559 1982 8615
rect 1842 2295 1898 2351
rect 1498 1908 1554 1964
rect 1498 864 1554 920
rect 2178 3491 2234 3547
rect 2094 1543 2150 1599
rect 4326 11338 4382 11340
rect 4326 11286 4328 11338
rect 4328 11286 4380 11338
rect 4380 11286 4382 11338
rect 4326 11284 4382 11286
rect 4326 9924 4382 9926
rect 4326 9872 4328 9924
rect 4328 9872 4380 9924
rect 4380 9872 4382 9924
rect 4326 9870 4382 9872
rect 2864 8559 2920 8615
rect 4326 8510 4382 8512
rect 4326 8458 4328 8510
rect 4328 8458 4380 8510
rect 4380 8458 4382 8510
rect 4326 8456 4382 8458
rect 4326 7096 4382 7098
rect 4326 7044 4328 7096
rect 4328 7044 4380 7096
rect 4380 7044 4382 7096
rect 4326 7042 4382 7044
rect 4326 5682 4382 5684
rect 4326 5630 4328 5682
rect 4328 5630 4380 5682
rect 4380 5630 4382 5682
rect 4326 5628 4382 5630
rect 4326 4268 4382 4270
rect 4326 4216 4328 4268
rect 4328 4216 4380 4268
rect 4380 4216 4382 4268
rect 4326 4214 4382 4216
rect 3242 3545 3298 3547
rect 3242 3493 3244 3545
rect 3244 3493 3296 3545
rect 3296 3493 3298 3545
rect 3242 3491 3298 3493
rect 2346 2295 2402 2351
rect 2262 1908 2318 1964
rect 4326 2854 4382 2856
rect 4326 2802 4328 2854
rect 4328 2802 4380 2854
rect 4380 2802 4382 2854
rect 4326 2800 4382 2802
rect 2514 2282 2570 2338
rect 3265 2336 3321 2338
rect 3265 2284 3267 2336
rect 3267 2284 3319 2336
rect 3319 2284 3321 2336
rect 3265 2282 3321 2284
rect 3610 1543 3666 1599
rect 4326 1440 4382 1442
rect 4326 1388 4328 1440
rect 4328 1388 4380 1440
rect 4380 1388 4382 1440
rect 4326 1386 4382 1388
rect 2514 864 2570 920
rect 2430 113 2486 169
rect 4264 113 4320 169
rect 4326 26 4382 28
rect 4326 -26 4328 26
rect 4328 -26 4380 26
rect 4380 -26 4382 26
rect 4326 -28 4382 -26
<< metal3 >>
rect 399 21503 497 21601
rect 1135 21503 1233 21601
rect 399 20383 497 20481
rect 1135 20383 1233 20481
rect 399 19263 497 19361
rect 1135 19263 1233 19361
rect 399 18143 497 18241
rect 1135 18143 1233 18241
rect 399 17023 497 17121
rect 1135 17023 1233 17121
rect 399 15903 497 16001
rect 1135 15903 1233 16001
rect 399 14783 497 14881
rect 1135 14783 1233 14881
rect 399 13663 497 13761
rect 1135 13663 1233 13761
rect 399 12543 497 12641
rect 1135 12543 1233 12641
rect 399 11423 497 11521
rect 1135 11423 1233 11521
rect 4305 11340 4403 11361
rect 4305 11284 4326 11340
rect 4382 11284 4403 11340
rect 4305 11263 4403 11284
rect 4305 9926 4403 9947
rect 4305 9870 4326 9926
rect 4382 9870 4403 9926
rect 4305 9849 4403 9870
rect 1921 8617 1987 8620
rect 2859 8617 2925 8620
rect 1921 8615 2925 8617
rect 1921 8559 1926 8615
rect 1982 8559 2864 8615
rect 2920 8559 2925 8615
rect 1921 8557 2925 8559
rect 1921 8554 1987 8557
rect 2859 8554 2925 8557
rect 4305 8512 4403 8533
rect 4305 8456 4326 8512
rect 4382 8456 4403 8512
rect 4305 8435 4403 8456
rect 4305 7098 4403 7119
rect 4305 7042 4326 7098
rect 4382 7042 4403 7098
rect 4305 7021 4403 7042
rect 4305 5684 4403 5705
rect 4305 5628 4326 5684
rect 4382 5628 4403 5684
rect 4305 5607 4403 5628
rect 4305 4270 4403 4291
rect 4305 4214 4326 4270
rect 4382 4214 4403 4270
rect 4305 4193 4403 4214
rect 2173 3549 2239 3552
rect 3237 3549 3303 3552
rect 2173 3547 3303 3549
rect 2173 3491 2178 3547
rect 2234 3491 3242 3547
rect 3298 3491 3303 3547
rect 2173 3489 3303 3491
rect 2173 3486 2239 3489
rect 3237 3486 3303 3489
rect -49 2781 49 2879
rect 4305 2856 4403 2877
rect 4305 2800 4326 2856
rect 4382 2800 4403 2856
rect 4305 2779 4403 2800
rect 1837 2353 1903 2356
rect 2341 2353 2407 2356
rect 1837 2351 2407 2353
rect 1837 2295 1842 2351
rect 1898 2295 2346 2351
rect 2402 2295 2407 2351
rect 1837 2293 2407 2295
rect 1837 2290 1903 2293
rect 2341 2290 2407 2293
rect 2509 2340 2575 2343
rect 3260 2340 3326 2343
rect 2509 2338 3326 2340
rect 2509 2282 2514 2338
rect 2570 2282 3265 2338
rect 3321 2282 3326 2338
rect 2509 2280 3326 2282
rect 2509 2277 2575 2280
rect 3260 2277 3326 2280
rect 1493 1966 1559 1969
rect 2257 1966 2323 1969
rect 1493 1964 2323 1966
rect 1493 1908 1498 1964
rect 1554 1908 2262 1964
rect 2318 1908 2323 1964
rect 1493 1906 2323 1908
rect 1493 1903 1559 1906
rect 2257 1903 2323 1906
rect 2089 1601 2155 1604
rect 3605 1601 3671 1604
rect 2089 1599 3671 1601
rect 2089 1543 2094 1599
rect 2150 1543 3610 1599
rect 3666 1543 3671 1599
rect 2089 1541 3671 1543
rect 2089 1538 2155 1541
rect 3605 1538 3671 1541
rect -49 1365 49 1463
rect 4305 1442 4403 1463
rect 4305 1386 4326 1442
rect 4382 1386 4403 1442
rect 4305 1365 4403 1386
rect 1493 922 1559 925
rect 2509 922 2575 925
rect 1493 920 2575 922
rect 1493 864 1498 920
rect 1554 864 2514 920
rect 2570 864 2575 920
rect 1493 862 2575 864
rect 1493 859 1559 862
rect 2509 859 2575 862
rect 2425 171 2491 174
rect 4259 171 4325 174
rect 2425 169 4325 171
rect 2425 113 2430 169
rect 2486 113 4264 169
rect 4320 113 4325 169
rect 2425 111 4325 113
rect 2425 108 2491 111
rect 4259 108 4325 111
rect -49 -51 49 47
rect 4305 28 4403 33
rect 4305 -28 4326 28
rect 4382 -28 4403 28
rect 4305 -49 4403 -28
use contact_32  contact_32_9
timestamp 1636140361
transform 1 0 1921 0 1 8550
box 0 0 1 1
use contact_8  contact_8_26
timestamp 1636140361
transform 1 0 1922 0 1 6018
box 0 0 1 1
use contact_8  contact_8_24
timestamp 1636140361
transform 1 0 171 0 1 7021
box 0 0 1 1
use contact_9  contact_9_12
timestamp 1636140361
transform 1 0 1837 0 1 2286
box 0 0 1 1
use contact_8  contact_8_21
timestamp 1636140361
transform 1 0 351 0 1 4210
box 0 0 1 1
use dff_buf_array  dff_buf_array_0
timestamp 1636140361
transform 1 0 0 0 1 0
box -49 -51 1976 2879
use contact_9  contact_9_11
timestamp 1636140361
transform 1 0 1493 0 1 855
box 0 0 1 1
use contact_9  contact_9_10
timestamp 1636140361
transform 1 0 1493 0 1 1899
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1636140361
transform 1 0 2748 0 1 636
box 0 0 1 1
use pinv_0  pinv_0_0
timestamp 1636140361
transform 1 0 2696 0 -1 2828
box -36 -17 404 1471
use contact_32  contact_32_3
timestamp 1636140361
transform 1 0 2509 0 1 855
box 0 0 1 1
use contact_32  contact_32_6
timestamp 1636140361
transform 1 0 2425 0 1 104
box 0 0 1 1
use contact_8  contact_8_14
timestamp 1636140361
transform 1 0 2745 0 1 637
box 0 0 1 1
use pand2_0  pand2_0_1
timestamp 1636140361
transform 1 0 3064 0 -1 2828
box -36 -17 782 1471
use pdriver_1  pdriver_1_0
timestamp 1636140361
transform 1 0 2696 0 1 0
box -36 -17 1694 1471
use contact_32  contact_32_8
timestamp 1636140361
transform 1 0 2089 0 1 1534
box 0 0 1 1
use pand2_0  pand2_0_0
timestamp 1636140361
transform 1 0 2696 0 1 2828
box -36 -17 782 1471
use contact_8  contact_8_13
timestamp 1636140361
transform 1 0 2426 0 1 2127
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1636140361
transform 1 0 2748 0 1 2126
box 0 0 1 1
use contact_32  contact_32_5
timestamp 1636140361
transform 1 0 2509 0 1 2273
box 0 0 1 1
use contact_32  contact_32_4
timestamp 1636140361
transform 1 0 2257 0 1 1899
box 0 0 1 1
use contact_32  contact_32_2
timestamp 1636140361
transform 1 0 2341 0 1 2286
box 0 0 1 1
use contact_7  contact_7_19
timestamp 1636140361
transform 1 0 3264 0 1 2277
box 0 0 1 1
use contact_8  contact_8_19
timestamp 1636140361
transform 1 0 3261 0 1 2278
box 0 0 1 1
use contact_9  contact_9_9
timestamp 1636140361
transform 1 0 3260 0 1 2273
box 0 0 1 1
use contact_7  contact_7_18
timestamp 1636140361
transform 1 0 3264 0 1 2277
box 0 0 1 1
use contact_8  contact_8_18
timestamp 1636140361
transform 1 0 3261 0 1 2278
box 0 0 1 1
use contact_9  contact_9_8
timestamp 1636140361
transform 1 0 3260 0 1 2273
box 0 0 1 1
use contact_32  contact_32_1
timestamp 1636140361
transform 1 0 3605 0 1 1534
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1636140361
transform 1 0 3609 0 1 2104
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1636140361
transform 1 0 3606 0 1 2105
box 0 0 1 1
use contact_32  contact_32_7
timestamp 1636140361
transform 1 0 2173 0 1 3482
box 0 0 1 1
use contact_8  contact_8_11
timestamp 1636140361
transform 1 0 2426 0 1 3066
box 0 0 1 1
use contact_8  contact_8_15
timestamp 1636140361
transform 1 0 2510 0 1 3314
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1636140361
transform 1 0 2896 0 1 3313
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1636140361
transform 1 0 2796 0 1 3065
box 0 0 1 1
use contact_8  contact_8_16
timestamp 1636140361
transform 1 0 3238 0 1 3487
box 0 0 1 1
use contact_7  contact_7_16
timestamp 1636140361
transform 1 0 3241 0 1 3486
box 0 0 1 1
use contact_9  contact_9_7
timestamp 1636140361
transform 1 0 3237 0 1 3482
box 0 0 1 1
use contact_8  contact_8_17
timestamp 1636140361
transform 1 0 3238 0 1 3487
box 0 0 1 1
use contact_7  contact_7_17
timestamp 1636140361
transform 1 0 3241 0 1 3486
box 0 0 1 1
use contact_8  contact_8_12
timestamp 1636140361
transform 1 0 2426 0 1 4210
box 0 0 1 1
use pdriver_2  pdriver_2_0
timestamp 1636140361
transform 1 0 2696 0 -1 5656
box -36 -17 1694 1471
use contact_7  contact_7_11
timestamp 1636140361
transform 1 0 2748 0 1 4954
box 0 0 1 1
use contact_8  contact_8_20
timestamp 1636140361
transform 1 0 2090 0 1 4955
box 0 0 1 1
use contact_7  contact_7_25
timestamp 1636140361
transform 1 0 2763 0 1 5893
box 0 0 1 1
use contact_8  contact_8_30
timestamp 1636140361
transform 1 0 2258 0 1 5894
box 0 0 1 1
use pand3  pand3_0
timestamp 1636140361
transform 1 0 2696 0 1 5656
box -36 -17 882 1471
use contact_8  contact_8_23
timestamp 1636140361
transform 1 0 2006 0 1 7021
box 0 0 1 1
use contact_8  contact_8_25
timestamp 1636140361
transform 1 0 2090 0 1 6142
box 0 0 1 1
use contact_7  contact_7_21
timestamp 1636140361
transform 1 0 3029 0 1 6141
box 0 0 1 1
use contact_7  contact_7_24
timestamp 1636140361
transform 1 0 2896 0 1 6017
box 0 0 1 1
use pnand2_1  pnand2_1_0
timestamp 1636140361
transform 1 0 2696 0 -1 8484
box -36 -17 504 1471
use contact_8  contact_8_39
timestamp 1636140361
transform 1 0 3338 0 1 6331
box 0 0 1 1
use contact_7  contact_7_37
timestamp 1636140361
transform 1 0 3341 0 1 6330
box 0 0 1 1
use pdriver_5  pdriver_5_0
timestamp 1636140361
transform 1 0 3164 0 -1 8484
box -36 -17 1178 1471
use contact_8  contact_8_22
timestamp 1636140361
transform 1 0 2006 0 1 7934
box 0 0 1 1
use contact_32  contact_32_10
timestamp 1636140361
transform 1 0 2859 0 1 8550
box 0 0 1 1
use contact_7  contact_7_20
timestamp 1636140361
transform 1 0 2896 0 1 7933
box 0 0 1 1
use contact_7  contact_7_22
timestamp 1636140361
transform 1 0 2796 0 1 8181
box 0 0 1 1
use contact_8  contact_8_29
timestamp 1636140361
transform 1 0 2174 0 1 8182
box 0 0 1 1
use pinv_0  pinv_0_1
timestamp 1636140361
transform 1 0 2696 0 1 8484
box -36 -17 404 1471
use contact_8  contact_8_27
timestamp 1636140361
transform 1 0 2006 0 1 9121
box 0 0 1 1
use contact_8  contact_8_28
timestamp 1636140361
transform 1 0 2860 0 1 9121
box 0 0 1 1
use contact_7  contact_7_23
timestamp 1636140361
transform 1 0 2863 0 1 9120
box 0 0 1 1
use contact_7  contact_7_26
timestamp 1636140361
transform 1 0 2748 0 1 9120
box 0 0 1 1
use pand3_0  pand3_0_0
timestamp 1636140361
transform 1 0 2696 0 -1 11312
box -36 -17 882 1471
use contact_9  contact_9_3
timestamp 1636140361
transform 1 0 4321 0 1 -37
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1636140361
transform 1 0 4322 0 1 -32
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1636140361
transform 1 0 4325 0 1 -33
box 0 0 1 1
use contact_32  contact_32_0
timestamp 1636140361
transform 1 0 4259 0 1 104
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1636140361
transform 1 0 4263 0 1 674
box 0 0 1 1
use contact_8  contact_8_8
timestamp 1636140361
transform 1 0 4260 0 1 675
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1636140361
transform 1 0 4263 0 1 674
box 0 0 1 1
use contact_8  contact_8_9
timestamp 1636140361
transform 1 0 4260 0 1 675
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1636140361
transform 1 0 4321 0 1 1377
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1636140361
transform 1 0 4322 0 1 1382
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1636140361
transform 1 0 4325 0 1 1381
box 0 0 1 1
use contact_9  contact_9_4
timestamp 1636140361
transform 1 0 4321 0 1 1377
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1636140361
transform 1 0 4322 0 1 1382
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1636140361
transform 1 0 4325 0 1 1381
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1636140361
transform 1 0 4322 0 1 2796
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1636140361
transform 1 0 4325 0 1 2795
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1636140361
transform 1 0 4321 0 1 2791
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1636140361
transform 1 0 4322 0 1 2796
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1636140361
transform 1 0 4325 0 1 2795
box 0 0 1 1
use contact_9  contact_9_6
timestamp 1636140361
transform 1 0 4321 0 1 2791
box 0 0 1 1
use contact_9  contact_9_0
timestamp 1636140361
transform 1 0 4321 0 1 4205
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1636140361
transform 1 0 4322 0 1 4210
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1636140361
transform 1 0 4325 0 1 4209
box 0 0 1 1
use contact_9  contact_9_5
timestamp 1636140361
transform 1 0 4321 0 1 4205
box 0 0 1 1
use contact_8  contact_8_10
timestamp 1636140361
transform 1 0 4322 0 1 4210
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1636140361
transform 1 0 4325 0 1 4209
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1636140361
transform 1 0 4260 0 1 4917
box 0 0 1 1
use contact_7  contact_7_0
timestamp 1636140361
transform 1 0 4263 0 1 4916
box 0 0 1 1
use contact_9  contact_9_18
timestamp 1636140361
transform 1 0 4321 0 1 5619
box 0 0 1 1
use contact_8  contact_8_36
timestamp 1636140361
transform 1 0 4322 0 1 5624
box 0 0 1 1
use contact_7  contact_7_32
timestamp 1636140361
transform 1 0 4325 0 1 5623
box 0 0 1 1
use contact_9  contact_9_20
timestamp 1636140361
transform 1 0 4321 0 1 5619
box 0 0 1 1
use contact_8  contact_8_38
timestamp 1636140361
transform 1 0 4322 0 1 5624
box 0 0 1 1
use contact_7  contact_7_34
timestamp 1636140361
transform 1 0 4325 0 1 5623
box 0 0 1 1
use contact_9  contact_9_17
timestamp 1636140361
transform 1 0 4321 0 1 7033
box 0 0 1 1
use contact_8  contact_8_35
timestamp 1636140361
transform 1 0 4322 0 1 7038
box 0 0 1 1
use contact_7  contact_7_31
timestamp 1636140361
transform 1 0 4325 0 1 7037
box 0 0 1 1
use contact_9  contact_9_19
timestamp 1636140361
transform 1 0 4321 0 1 7033
box 0 0 1 1
use contact_8  contact_8_37
timestamp 1636140361
transform 1 0 4322 0 1 7038
box 0 0 1 1
use contact_7  contact_7_33
timestamp 1636140361
transform 1 0 4325 0 1 7037
box 0 0 1 1
use contact_7  contact_7_35
timestamp 1636140361
transform 1 0 4215 0 1 7744
box 0 0 1 1
use contact_8  contact_8_41
timestamp 1636140361
transform 1 0 4212 0 1 7745
box 0 0 1 1
use contact_9  contact_9_14
timestamp 1636140361
transform 1 0 4321 0 1 8447
box 0 0 1 1
use contact_8  contact_8_32
timestamp 1636140361
transform 1 0 4322 0 1 8452
box 0 0 1 1
use contact_7  contact_7_28
timestamp 1636140361
transform 1 0 4325 0 1 8451
box 0 0 1 1
use contact_9  contact_9_16
timestamp 1636140361
transform 1 0 4321 0 1 8447
box 0 0 1 1
use contact_8  contact_8_34
timestamp 1636140361
transform 1 0 4322 0 1 8452
box 0 0 1 1
use contact_7  contact_7_30
timestamp 1636140361
transform 1 0 4325 0 1 8451
box 0 0 1 1
use contact_9  contact_9_13
timestamp 1636140361
transform 1 0 4321 0 1 9861
box 0 0 1 1
use contact_8  contact_8_31
timestamp 1636140361
transform 1 0 4322 0 1 9866
box 0 0 1 1
use contact_7  contact_7_27
timestamp 1636140361
transform 1 0 4325 0 1 9865
box 0 0 1 1
use contact_9  contact_9_15
timestamp 1636140361
transform 1 0 4321 0 1 9861
box 0 0 1 1
use contact_8  contact_8_33
timestamp 1636140361
transform 1 0 4322 0 1 9866
box 0 0 1 1
use contact_7  contact_7_29
timestamp 1636140361
transform 1 0 4325 0 1 9865
box 0 0 1 1
use delay_chain  delay_chain_0
timestamp 1636140361
transform -1 0 1840 0 1 11472
box -36 -49 1876 10137
use contact_8  contact_8_45
timestamp 1636140361
transform 1 0 2342 0 1 10762
box 0 0 1 1
use contact_7  contact_7_41
timestamp 1636140361
transform 1 0 3029 0 1 10761
box 0 0 1 1
use contact_7  contact_7_40
timestamp 1636140361
transform 1 0 2763 0 1 11009
box 0 0 1 1
use contact_7  contact_7_39
timestamp 1636140361
transform 1 0 2896 0 1 10885
box 0 0 1 1
use contact_8  contact_8_43
timestamp 1636140361
transform 1 0 2006 0 1 11010
box 0 0 1 1
use contact_8  contact_8_42
timestamp 1636140361
transform 1 0 2090 0 1 10886
box 0 0 1 1
use contact_7  contact_7_36
timestamp 1636140361
transform 1 0 3341 0 1 10572
box 0 0 1 1
use contact_8  contact_8_40
timestamp 1636140361
transform 1 0 3338 0 1 10573
box 0 0 1 1
use contact_7  contact_7_38
timestamp 1636140361
transform 1 0 4325 0 1 11279
box 0 0 1 1
use contact_8  contact_8_44
timestamp 1636140361
transform 1 0 4322 0 1 11280
box 0 0 1 1
use contact_9  contact_9_21
timestamp 1636140361
transform 1 0 4321 0 1 11275
box 0 0 1 1
<< labels >>
rlabel metal2 s 1762 11733 1762 11733 4 rbl_bl
port 4 nsew
rlabel metal2 s 4341 7777 4341 7777 4 p_en_bar
port 7 nsew
rlabel metal2 s 170 564 170 564 4 csb
port 1 nsew
rlabel metal2 s 3904 6363 3904 6363 4 w_en
port 6 nsew
rlabel metal2 s 3904 10605 3904 10605 4 s_en
port 5 nsew
rlabel metal2 s 4365 707 4365 707 4 clk_buf
port 9 nsew
rlabel metal2 s 2777 669 2777 669 4 clk
port 3 nsew
rlabel metal2 s 170 2264 170 2264 4 web
port 2 nsew
rlabel metal2 s 4365 4949 4365 4949 4 wl_en
port 8 nsew
rlabel metal3 s 448 12592 448 12592 4 vdd
port 10 nsew
rlabel metal3 s 1184 17072 1184 17072 4 vdd
port 10 nsew
rlabel metal3 s 448 14832 448 14832 4 vdd
port 10 nsew
rlabel metal3 s 448 19312 448 19312 4 vdd
port 10 nsew
rlabel metal3 s 448 21552 448 21552 4 vdd
port 10 nsew
rlabel metal3 s 1184 14832 1184 14832 4 vdd
port 10 nsew
rlabel metal3 s 1184 21552 1184 21552 4 vdd
port 10 nsew
rlabel metal3 s 4354 9898 4354 9898 4 vdd
port 10 nsew
rlabel metal3 s 1184 12592 1184 12592 4 vdd
port 10 nsew
rlabel metal3 s 448 17072 448 17072 4 vdd
port 10 nsew
rlabel metal3 s 0 1414 0 1414 4 vdd
port 10 nsew
rlabel metal3 s 4354 4242 4354 4242 4 vdd
port 10 nsew
rlabel metal3 s 1184 19312 1184 19312 4 vdd
port 10 nsew
rlabel metal3 s 4354 1414 4354 1414 4 vdd
port 10 nsew
rlabel metal3 s 4354 7070 4354 7070 4 vdd
port 10 nsew
rlabel metal3 s 4354 11312 4354 11312 4 gnd
port 11 nsew
rlabel metal3 s 4354 8484 4354 8484 4 gnd
port 11 nsew
rlabel metal3 s 1184 11472 1184 11472 4 gnd
port 11 nsew
rlabel metal3 s 1184 18192 1184 18192 4 gnd
port 11 nsew
rlabel metal3 s 1184 20432 1184 20432 4 gnd
port 11 nsew
rlabel metal3 s 0 -2 0 -2 4 gnd
port 11 nsew
rlabel metal3 s 1184 13712 1184 13712 4 gnd
port 11 nsew
rlabel metal3 s 1184 15952 1184 15952 4 gnd
port 11 nsew
rlabel metal3 s 448 20432 448 20432 4 gnd
port 11 nsew
rlabel metal3 s 448 15952 448 15952 4 gnd
port 11 nsew
rlabel metal3 s 448 18192 448 18192 4 gnd
port 11 nsew
rlabel metal3 s 4354 0 4354 0 4 gnd
port 11 nsew
rlabel metal3 s 448 13712 448 13712 4 gnd
port 11 nsew
rlabel metal3 s 4354 2828 4354 2828 4 gnd
port 11 nsew
rlabel metal3 s 0 2830 0 2830 4 gnd
port 11 nsew
rlabel metal3 s 4354 5656 4354 5656 4 gnd
port 11 nsew
rlabel metal3 s 448 11472 448 11472 4 gnd
port 11 nsew
<< properties >>
string FIXED_BBOX 4321 -37 4387 0
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_END 6443502
string GDS_START 6425666
<< end >>
