magic
tech sky130A
magscale 1 2
timestamp 1636140361
<< checkpaint >>
rect -1296 -1277 3500 2731
<< nwell >>
rect -36 679 2240 1471
<< pwell >>
rect 2068 25 2170 159
<< psubdiff >>
rect 2094 109 2144 133
rect 2094 75 2102 109
rect 2136 75 2144 109
rect 2094 51 2144 75
<< nsubdiff >>
rect 2094 1339 2144 1363
rect 2094 1305 2102 1339
rect 2136 1305 2144 1339
rect 2094 1281 2144 1305
<< psubdiffcont >>
rect 2102 75 2136 109
<< nsubdiffcont >>
rect 2102 1305 2136 1339
<< poly >>
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 2204 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 1138 1130 1172 1397
rect 1354 1130 1388 1397
rect 1570 1130 1604 1397
rect 1786 1130 1820 1397
rect 1998 1130 2032 1397
rect 2102 1339 2136 1397
rect 2102 1289 2136 1305
rect 64 724 98 740
rect 64 674 98 690
rect 1030 724 1064 1096
rect 1030 690 1081 724
rect 1030 318 1064 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 1138 17 1172 218
rect 1354 17 1388 218
rect 1570 17 1604 218
rect 1786 17 1820 218
rect 1998 17 2032 218
rect 2102 109 2136 125
rect 2102 17 2136 75
rect 0 -17 2204 17
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_16  sky130_sram_1kbyte_1rw1r_32x256_8_contact_16_0
timestamp 1636140361
transform 1 0 48 0 1 674
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_29  sky130_sram_1kbyte_1rw1r_32x256_8_contact_29_0
timestamp 1636140361
transform 1 0 2094 0 1 51
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_28  sky130_sram_1kbyte_1rw1r_32x256_8_contact_28_0
timestamp 1636140361
transform 1 0 2094 0 1 1281
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m18_w2_000_sli_dli_da_p  sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m18_w2_000_sli_dli_da_p_0
timestamp 1636140361
transform 1 0 54 0 1 51
box -26 -26 2012 456
use sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m18_w2_000_sli_dli_da_p  sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m18_w2_000_sli_dli_da_p_0
timestamp 1636140361
transform 1 0 54 0 1 963
box -59 -56 2045 454
<< labels >>
rlabel locali s 81 707 81 707 4 A
port 1 nsew
rlabel locali s 1064 707 1064 707 4 Z
port 2 nsew
rlabel locali s 1102 0 1102 0 4 gnd
port 3 nsew
rlabel locali s 1102 1414 1102 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2204 1414
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_END 100586
string GDS_START 97564
<< end >>
