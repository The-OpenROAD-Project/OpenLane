magic
tech sky130A
magscale 1 2
timestamp 1636140361
<< checkpaint >>
rect 4284 -4490 50221 5721
<< metal1 >>
rect 13910 4398 13916 4450
rect 13968 4398 13974 4450
rect 18902 4398 18908 4450
rect 18960 4398 18966 4450
rect 23894 4398 23900 4450
rect 23952 4398 23958 4450
rect 28886 4398 28892 4450
rect 28944 4398 28950 4450
rect 33878 4398 33884 4450
rect 33936 4398 33942 4450
rect 38870 4398 38876 4450
rect 38928 4398 38934 4450
rect 43862 4398 43868 4450
rect 43920 4398 43926 4450
rect 48854 4398 48860 4450
rect 48912 4398 48918 4450
<< via1 >>
rect 13916 4398 13968 4450
rect 18908 4398 18960 4450
rect 23900 4398 23952 4450
rect 28892 4398 28944 4450
rect 33884 4398 33936 4450
rect 38876 4398 38928 4450
rect 43868 4398 43920 4450
rect 48860 4398 48912 4450
<< metal2 >>
rect 13914 4452 13970 4461
rect 13914 4387 13970 4396
rect 18906 4452 18962 4461
rect 18906 4387 18962 4396
rect 23898 4452 23954 4461
rect 23898 4387 23954 4396
rect 28890 4452 28946 4461
rect 28890 4387 28946 4396
rect 33882 4452 33938 4461
rect 33882 4387 33938 4396
rect 38874 4452 38930 4461
rect 38874 4387 38930 4396
rect 43866 4452 43922 4461
rect 43866 4387 43922 4396
rect 48858 4452 48914 4461
rect 48858 4387 48914 4396
rect 13629 3332 13685 3341
rect 13629 3267 13685 3276
rect 5591 -3165 5647 -3156
rect 5591 -3230 5647 -3221
rect 6759 -3165 6815 -3156
rect 6759 -3230 6815 -3221
rect 7927 -3165 7983 -3156
rect 7927 -3230 7983 -3221
rect 9095 -3165 9151 -3156
rect 9095 -3230 9151 -3221
rect 10263 -3165 10319 -3156
rect 10263 -3230 10319 -3221
rect 11431 -3165 11487 -3156
rect 11431 -3230 11487 -3221
rect 12599 -3165 12655 -3156
rect 12599 -3230 12655 -3221
rect 13767 -3165 13823 -3156
rect 13767 -3230 13823 -3221
rect 14935 -3165 14991 -3156
rect 14935 -3230 14991 -3221
<< via2 >>
rect 13914 4450 13970 4452
rect 13914 4398 13916 4450
rect 13916 4398 13968 4450
rect 13968 4398 13970 4450
rect 13914 4396 13970 4398
rect 18906 4450 18962 4452
rect 18906 4398 18908 4450
rect 18908 4398 18960 4450
rect 18960 4398 18962 4450
rect 18906 4396 18962 4398
rect 23898 4450 23954 4452
rect 23898 4398 23900 4450
rect 23900 4398 23952 4450
rect 23952 4398 23954 4450
rect 23898 4396 23954 4398
rect 28890 4450 28946 4452
rect 28890 4398 28892 4450
rect 28892 4398 28944 4450
rect 28944 4398 28946 4450
rect 28890 4396 28946 4398
rect 33882 4450 33938 4452
rect 33882 4398 33884 4450
rect 33884 4398 33936 4450
rect 33936 4398 33938 4450
rect 33882 4396 33938 4398
rect 38874 4450 38930 4452
rect 38874 4398 38876 4450
rect 38876 4398 38928 4450
rect 38928 4398 38930 4450
rect 38874 4396 38930 4398
rect 43866 4450 43922 4452
rect 43866 4398 43868 4450
rect 43868 4398 43920 4450
rect 43920 4398 43922 4450
rect 43866 4396 43922 4398
rect 48858 4450 48914 4452
rect 48858 4398 48860 4450
rect 48860 4398 48912 4450
rect 48912 4398 48914 4450
rect 48858 4396 48914 4398
rect 13629 3276 13685 3332
rect 5591 -3221 5647 -3165
rect 6759 -3221 6815 -3165
rect 7927 -3221 7983 -3165
rect 9095 -3221 9151 -3165
rect 10263 -3221 10319 -3165
rect 11431 -3221 11487 -3165
rect 12599 -3221 12655 -3165
rect 13767 -3221 13823 -3165
rect 14935 -3221 14991 -3165
<< metal3 >>
rect 13909 4456 13975 4457
rect 18901 4456 18967 4457
rect 23893 4456 23959 4457
rect 28885 4456 28951 4457
rect 33877 4456 33943 4457
rect 38869 4456 38935 4457
rect 43861 4456 43927 4457
rect 48853 4456 48919 4457
rect 13867 4392 13910 4456
rect 13974 4392 14017 4456
rect 18859 4392 18902 4456
rect 18966 4392 19009 4456
rect 23851 4392 23894 4456
rect 23958 4392 24001 4456
rect 28843 4392 28886 4456
rect 28950 4392 28993 4456
rect 33835 4392 33878 4456
rect 33942 4392 33985 4456
rect 38827 4392 38870 4456
rect 38934 4392 38977 4456
rect 43819 4392 43862 4456
rect 43926 4392 43969 4456
rect 48811 4392 48854 4456
rect 48918 4392 48961 4456
rect 13909 4391 13975 4392
rect 18901 4391 18967 4392
rect 23893 4391 23959 4392
rect 28885 4391 28951 4392
rect 33877 4391 33943 4392
rect 38869 4391 38935 4392
rect 43861 4391 43927 4392
rect 48853 4391 48919 4392
rect 13624 3336 13690 3337
rect 13582 3272 13625 3336
rect 13689 3272 13732 3336
rect 13624 3271 13690 3272
rect 6749 -516 6755 -452
rect 6819 -454 6825 -452
rect 13904 -454 13910 -452
rect 6819 -514 13910 -454
rect 6819 -516 6825 -514
rect 13904 -516 13910 -514
rect 13974 -516 13980 -452
rect 5581 -760 5587 -696
rect 5651 -698 5657 -696
rect 13619 -698 13625 -696
rect 5651 -758 13625 -698
rect 5651 -760 5657 -758
rect 13619 -760 13625 -758
rect 13689 -760 13695 -696
rect 14925 -760 14931 -696
rect 14995 -698 15001 -696
rect 48848 -698 48854 -696
rect 14995 -758 48854 -698
rect 14995 -760 15001 -758
rect 48848 -760 48854 -758
rect 48918 -760 48924 -696
rect 13757 -1004 13763 -940
rect 13827 -942 13833 -940
rect 43856 -942 43862 -940
rect 13827 -1002 43862 -942
rect 13827 -1004 13833 -1002
rect 43856 -1004 43862 -1002
rect 43926 -1004 43932 -940
rect 12589 -1248 12595 -1184
rect 12659 -1186 12665 -1184
rect 38864 -1186 38870 -1184
rect 12659 -1246 38870 -1186
rect 12659 -1248 12665 -1246
rect 38864 -1248 38870 -1246
rect 38934 -1248 38940 -1184
rect 11421 -1492 11427 -1428
rect 11491 -1430 11497 -1428
rect 33872 -1430 33878 -1428
rect 11491 -1490 33878 -1430
rect 11491 -1492 11497 -1490
rect 33872 -1492 33878 -1490
rect 33942 -1492 33948 -1428
rect 10253 -1736 10259 -1672
rect 10323 -1674 10329 -1672
rect 28880 -1674 28886 -1672
rect 10323 -1734 28886 -1674
rect 10323 -1736 10329 -1734
rect 28880 -1736 28886 -1734
rect 28950 -1736 28956 -1672
rect 9085 -1980 9091 -1916
rect 9155 -1918 9161 -1916
rect 23888 -1918 23894 -1916
rect 9155 -1978 23894 -1918
rect 9155 -1980 9161 -1978
rect 23888 -1980 23894 -1978
rect 23958 -1980 23964 -1916
rect 7917 -2224 7923 -2160
rect 7987 -2162 7993 -2160
rect 18896 -2162 18902 -2160
rect 7987 -2222 18902 -2162
rect 7987 -2224 7993 -2222
rect 18896 -2224 18902 -2222
rect 18966 -2224 18972 -2160
rect 5586 -3161 5652 -3160
rect 6754 -3161 6820 -3160
rect 7922 -3161 7988 -3160
rect 9090 -3161 9156 -3160
rect 10258 -3161 10324 -3160
rect 11426 -3161 11492 -3160
rect 12594 -3161 12660 -3160
rect 13762 -3161 13828 -3160
rect 14930 -3161 14996 -3160
rect 5544 -3225 5587 -3161
rect 5651 -3225 5694 -3161
rect 6712 -3225 6755 -3161
rect 6819 -3225 6862 -3161
rect 7880 -3225 7923 -3161
rect 7987 -3225 8030 -3161
rect 9048 -3225 9091 -3161
rect 9155 -3225 9198 -3161
rect 10216 -3225 10259 -3161
rect 10323 -3225 10366 -3161
rect 11384 -3225 11427 -3161
rect 11491 -3225 11534 -3161
rect 12552 -3225 12595 -3161
rect 12659 -3225 12702 -3161
rect 13720 -3225 13763 -3161
rect 13827 -3225 13870 -3161
rect 14888 -3225 14931 -3161
rect 14995 -3225 15038 -3161
rect 5586 -3226 5652 -3225
rect 6754 -3226 6820 -3225
rect 7922 -3226 7988 -3225
rect 9090 -3226 9156 -3225
rect 10258 -3226 10324 -3225
rect 11426 -3226 11492 -3225
rect 12594 -3226 12660 -3225
rect 13762 -3226 13828 -3225
rect 14930 -3226 14996 -3225
<< via3 >>
rect 13910 4452 13974 4456
rect 13910 4396 13914 4452
rect 13914 4396 13970 4452
rect 13970 4396 13974 4452
rect 13910 4392 13974 4396
rect 18902 4452 18966 4456
rect 18902 4396 18906 4452
rect 18906 4396 18962 4452
rect 18962 4396 18966 4452
rect 18902 4392 18966 4396
rect 23894 4452 23958 4456
rect 23894 4396 23898 4452
rect 23898 4396 23954 4452
rect 23954 4396 23958 4452
rect 23894 4392 23958 4396
rect 28886 4452 28950 4456
rect 28886 4396 28890 4452
rect 28890 4396 28946 4452
rect 28946 4396 28950 4452
rect 28886 4392 28950 4396
rect 33878 4452 33942 4456
rect 33878 4396 33882 4452
rect 33882 4396 33938 4452
rect 33938 4396 33942 4452
rect 33878 4392 33942 4396
rect 38870 4452 38934 4456
rect 38870 4396 38874 4452
rect 38874 4396 38930 4452
rect 38930 4396 38934 4452
rect 38870 4392 38934 4396
rect 43862 4452 43926 4456
rect 43862 4396 43866 4452
rect 43866 4396 43922 4452
rect 43922 4396 43926 4452
rect 43862 4392 43926 4396
rect 48854 4452 48918 4456
rect 48854 4396 48858 4452
rect 48858 4396 48914 4452
rect 48914 4396 48918 4452
rect 48854 4392 48918 4396
rect 13625 3332 13689 3336
rect 13625 3276 13629 3332
rect 13629 3276 13685 3332
rect 13685 3276 13689 3332
rect 13625 3272 13689 3276
rect 6755 -516 6819 -452
rect 13910 -516 13974 -452
rect 5587 -760 5651 -696
rect 13625 -760 13689 -696
rect 14931 -760 14995 -696
rect 48854 -760 48918 -696
rect 13763 -1004 13827 -940
rect 43862 -1004 43926 -940
rect 12595 -1248 12659 -1184
rect 38870 -1248 38934 -1184
rect 11427 -1492 11491 -1428
rect 33878 -1492 33942 -1428
rect 10259 -1736 10323 -1672
rect 28886 -1736 28950 -1672
rect 9091 -1980 9155 -1916
rect 23894 -1980 23958 -1916
rect 7923 -2224 7987 -2160
rect 18902 -2224 18966 -2160
rect 5587 -3165 5651 -3161
rect 5587 -3221 5591 -3165
rect 5591 -3221 5647 -3165
rect 5647 -3221 5651 -3165
rect 5587 -3225 5651 -3221
rect 6755 -3165 6819 -3161
rect 6755 -3221 6759 -3165
rect 6759 -3221 6815 -3165
rect 6815 -3221 6819 -3165
rect 6755 -3225 6819 -3221
rect 7923 -3165 7987 -3161
rect 7923 -3221 7927 -3165
rect 7927 -3221 7983 -3165
rect 7983 -3221 7987 -3165
rect 7923 -3225 7987 -3221
rect 9091 -3165 9155 -3161
rect 9091 -3221 9095 -3165
rect 9095 -3221 9151 -3165
rect 9151 -3221 9155 -3165
rect 9091 -3225 9155 -3221
rect 10259 -3165 10323 -3161
rect 10259 -3221 10263 -3165
rect 10263 -3221 10319 -3165
rect 10319 -3221 10323 -3165
rect 10259 -3225 10323 -3221
rect 11427 -3165 11491 -3161
rect 11427 -3221 11431 -3165
rect 11431 -3221 11487 -3165
rect 11487 -3221 11491 -3165
rect 11427 -3225 11491 -3221
rect 12595 -3165 12659 -3161
rect 12595 -3221 12599 -3165
rect 12599 -3221 12655 -3165
rect 12655 -3221 12659 -3165
rect 12595 -3225 12659 -3221
rect 13763 -3165 13827 -3161
rect 13763 -3221 13767 -3165
rect 13767 -3221 13823 -3165
rect 13823 -3221 13827 -3165
rect 13763 -3225 13827 -3221
rect 14931 -3165 14995 -3161
rect 14931 -3221 14935 -3165
rect 14935 -3221 14991 -3165
rect 14991 -3221 14995 -3165
rect 14931 -3225 14995 -3221
<< metal4 >>
rect 13909 4456 13975 4457
rect 13909 4392 13910 4456
rect 13974 4392 13975 4456
rect 13909 4391 13975 4392
rect 18901 4456 18967 4457
rect 18901 4392 18902 4456
rect 18966 4392 18967 4456
rect 18901 4391 18967 4392
rect 23893 4456 23959 4457
rect 23893 4392 23894 4456
rect 23958 4392 23959 4456
rect 23893 4391 23959 4392
rect 28885 4456 28951 4457
rect 28885 4392 28886 4456
rect 28950 4392 28951 4456
rect 28885 4391 28951 4392
rect 33877 4456 33943 4457
rect 33877 4392 33878 4456
rect 33942 4392 33943 4456
rect 33877 4391 33943 4392
rect 38869 4456 38935 4457
rect 38869 4392 38870 4456
rect 38934 4392 38935 4456
rect 38869 4391 38935 4392
rect 43861 4456 43927 4457
rect 43861 4392 43862 4456
rect 43926 4392 43927 4456
rect 43861 4391 43927 4392
rect 48853 4456 48919 4457
rect 48853 4392 48854 4456
rect 48918 4392 48919 4456
rect 48853 4391 48919 4392
rect 13624 3336 13690 3337
rect 13624 3272 13625 3336
rect 13689 3272 13690 3336
rect 13624 3271 13690 3272
rect 6754 -452 6820 -451
rect 6754 -516 6755 -452
rect 6819 -516 6820 -452
rect 6754 -517 6820 -516
rect 5586 -696 5652 -695
rect 5586 -760 5587 -696
rect 5651 -760 5652 -696
rect 5586 -761 5652 -760
rect 5589 -3160 5649 -761
rect 6757 -3160 6817 -517
rect 13627 -695 13687 3271
rect 13912 -451 13972 4391
rect 13909 -452 13975 -451
rect 13909 -516 13910 -452
rect 13974 -516 13975 -452
rect 13909 -517 13975 -516
rect 13624 -696 13690 -695
rect 13624 -760 13625 -696
rect 13689 -760 13690 -696
rect 13624 -761 13690 -760
rect 14930 -696 14996 -695
rect 14930 -760 14931 -696
rect 14995 -760 14996 -696
rect 14930 -761 14996 -760
rect 13762 -940 13828 -939
rect 13762 -1004 13763 -940
rect 13827 -1004 13828 -940
rect 13762 -1005 13828 -1004
rect 12594 -1184 12660 -1183
rect 12594 -1248 12595 -1184
rect 12659 -1248 12660 -1184
rect 12594 -1249 12660 -1248
rect 11426 -1428 11492 -1427
rect 11426 -1492 11427 -1428
rect 11491 -1492 11492 -1428
rect 11426 -1493 11492 -1492
rect 10258 -1672 10324 -1671
rect 10258 -1736 10259 -1672
rect 10323 -1736 10324 -1672
rect 10258 -1737 10324 -1736
rect 9090 -1916 9156 -1915
rect 9090 -1980 9091 -1916
rect 9155 -1980 9156 -1916
rect 9090 -1981 9156 -1980
rect 7922 -2160 7988 -2159
rect 7922 -2224 7923 -2160
rect 7987 -2224 7988 -2160
rect 7922 -2225 7988 -2224
rect 7925 -3160 7985 -2225
rect 9093 -3160 9153 -1981
rect 10261 -3160 10321 -1737
rect 11429 -3160 11489 -1493
rect 12597 -3160 12657 -1249
rect 13765 -3160 13825 -1005
rect 14933 -3160 14993 -761
rect 18904 -2159 18964 4391
rect 23896 -1915 23956 4391
rect 28888 -1671 28948 4391
rect 33880 -1427 33940 4391
rect 38872 -1183 38932 4391
rect 43864 -939 43924 4391
rect 48856 -695 48916 4391
rect 48853 -696 48919 -695
rect 48853 -760 48854 -696
rect 48918 -760 48919 -696
rect 48853 -761 48919 -760
rect 43861 -940 43927 -939
rect 43861 -1004 43862 -940
rect 43926 -1004 43927 -940
rect 43861 -1005 43927 -1004
rect 38869 -1184 38935 -1183
rect 38869 -1248 38870 -1184
rect 38934 -1248 38935 -1184
rect 38869 -1249 38935 -1248
rect 33877 -1428 33943 -1427
rect 33877 -1492 33878 -1428
rect 33942 -1492 33943 -1428
rect 33877 -1493 33943 -1492
rect 28885 -1672 28951 -1671
rect 28885 -1736 28886 -1672
rect 28950 -1736 28951 -1672
rect 28885 -1737 28951 -1736
rect 23893 -1916 23959 -1915
rect 23893 -1980 23894 -1916
rect 23958 -1980 23959 -1916
rect 23893 -1981 23959 -1980
rect 18901 -2160 18967 -2159
rect 18901 -2224 18902 -2160
rect 18966 -2224 18967 -2160
rect 18901 -2225 18967 -2224
rect 5586 -3161 5652 -3160
rect 5586 -3225 5587 -3161
rect 5651 -3225 5652 -3161
rect 5586 -3226 5652 -3225
rect 6754 -3161 6820 -3160
rect 6754 -3225 6755 -3161
rect 6819 -3225 6820 -3161
rect 6754 -3226 6820 -3225
rect 7922 -3161 7988 -3160
rect 7922 -3225 7923 -3161
rect 7987 -3225 7988 -3161
rect 7922 -3226 7988 -3225
rect 9090 -3161 9156 -3160
rect 9090 -3225 9091 -3161
rect 9155 -3225 9156 -3161
rect 9090 -3226 9156 -3225
rect 10258 -3161 10324 -3160
rect 10258 -3225 10259 -3161
rect 10323 -3225 10324 -3161
rect 10258 -3226 10324 -3225
rect 11426 -3161 11492 -3160
rect 11426 -3225 11427 -3161
rect 11491 -3225 11492 -3161
rect 11426 -3226 11492 -3225
rect 12594 -3161 12660 -3160
rect 12594 -3225 12595 -3161
rect 12659 -3225 12660 -3161
rect 12594 -3226 12660 -3225
rect 13762 -3161 13828 -3160
rect 13762 -3225 13763 -3161
rect 13827 -3225 13828 -3161
rect 13762 -3226 13828 -3225
rect 14930 -3161 14996 -3160
rect 14930 -3225 14931 -3161
rect 14995 -3225 14996 -3161
rect 14930 -3226 14996 -3225
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_0
timestamp 1636140361
transform 1 0 6749 0 1 -3226
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_0
timestamp 1636140361
transform 1 0 6754 0 1 -3230
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1
timestamp 1636140361
transform 1 0 6749 0 1 -517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2
timestamp 1636140361
transform 1 0 13904 0 1 4391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_1
timestamp 1636140361
transform 1 0 13909 0 1 4387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_0
timestamp 1636140361
transform 1 0 13910 0 1 4392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_3
timestamp 1636140361
transform 1 0 13904 0 1 -517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_4
timestamp 1636140361
transform 1 0 14925 0 1 -3226
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_2
timestamp 1636140361
transform 1 0 14930 0 1 -3230
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_5
timestamp 1636140361
transform 1 0 14925 0 1 -761
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_6
timestamp 1636140361
transform 1 0 48848 0 1 4391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_3
timestamp 1636140361
transform 1 0 48853 0 1 4387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_1
timestamp 1636140361
transform 1 0 48854 0 1 4392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_7
timestamp 1636140361
transform 1 0 48848 0 1 -761
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_8
timestamp 1636140361
transform 1 0 5581 0 1 -3226
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_4
timestamp 1636140361
transform 1 0 5586 0 1 -3230
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_9
timestamp 1636140361
transform 1 0 5581 0 1 -761
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_10
timestamp 1636140361
transform 1 0 13619 0 1 3271
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_5
timestamp 1636140361
transform 1 0 13624 0 1 3267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_11
timestamp 1636140361
transform 1 0 13619 0 1 -761
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_12
timestamp 1636140361
transform 1 0 13757 0 1 -3226
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_6
timestamp 1636140361
transform 1 0 13762 0 1 -3230
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_13
timestamp 1636140361
transform 1 0 13757 0 1 -1005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_14
timestamp 1636140361
transform 1 0 43856 0 1 4391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_7
timestamp 1636140361
transform 1 0 43861 0 1 4387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_2
timestamp 1636140361
transform 1 0 43862 0 1 4392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_15
timestamp 1636140361
transform 1 0 43856 0 1 -1005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_16
timestamp 1636140361
transform 1 0 12589 0 1 -3226
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_8
timestamp 1636140361
transform 1 0 12594 0 1 -3230
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_17
timestamp 1636140361
transform 1 0 12589 0 1 -1249
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_18
timestamp 1636140361
transform 1 0 38864 0 1 4391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_9
timestamp 1636140361
transform 1 0 38869 0 1 4387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_3
timestamp 1636140361
transform 1 0 38870 0 1 4392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_19
timestamp 1636140361
transform 1 0 38864 0 1 -1249
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_20
timestamp 1636140361
transform 1 0 11421 0 1 -3226
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_10
timestamp 1636140361
transform 1 0 11426 0 1 -3230
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_21
timestamp 1636140361
transform 1 0 11421 0 1 -1493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_22
timestamp 1636140361
transform 1 0 33872 0 1 4391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_11
timestamp 1636140361
transform 1 0 33877 0 1 4387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_4
timestamp 1636140361
transform 1 0 33878 0 1 4392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_23
timestamp 1636140361
transform 1 0 33872 0 1 -1493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_24
timestamp 1636140361
transform 1 0 10253 0 1 -3226
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_12
timestamp 1636140361
transform 1 0 10258 0 1 -3230
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_25
timestamp 1636140361
transform 1 0 10253 0 1 -1737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_26
timestamp 1636140361
transform 1 0 28880 0 1 4391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_13
timestamp 1636140361
transform 1 0 28885 0 1 4387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_5
timestamp 1636140361
transform 1 0 28886 0 1 4392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_27
timestamp 1636140361
transform 1 0 28880 0 1 -1737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_28
timestamp 1636140361
transform 1 0 9085 0 1 -3226
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_14
timestamp 1636140361
transform 1 0 9090 0 1 -3230
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_29
timestamp 1636140361
transform 1 0 9085 0 1 -1981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_30
timestamp 1636140361
transform 1 0 23888 0 1 4391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_15
timestamp 1636140361
transform 1 0 23893 0 1 4387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_6
timestamp 1636140361
transform 1 0 23894 0 1 4392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_31
timestamp 1636140361
transform 1 0 23888 0 1 -1981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_32
timestamp 1636140361
transform 1 0 7917 0 1 -3226
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_16
timestamp 1636140361
transform 1 0 7922 0 1 -3230
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_33
timestamp 1636140361
transform 1 0 7917 0 1 -2225
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_34
timestamp 1636140361
transform 1 0 18896 0 1 4391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_17
timestamp 1636140361
transform 1 0 18901 0 1 4387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_7
timestamp 1636140361
transform 1 0 18902 0 1 4392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_35
timestamp 1636140361
transform 1 0 18896 0 1 -2225
box 0 0 1 1
<< properties >>
string FIXED_BBOX 5544 -3230 48961 4461
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_END 7031534
string GDS_START 7023422
<< end >>
