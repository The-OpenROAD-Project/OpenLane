VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS
MACRO digital_out_pad
   CLASS BLOCK ;
   FOREIGN digital_out_pad ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 80.0000 BY 165.0000 ;
   PIN in3v
      PORT
         LAYER met2 ;
	    RECT 63.940000 0.000000 64.980000 4.000000 ;
      END
   END in3v
   PIN in
      PORT
         LAYER met2 ;
	    RECT 65.970000 0.000000 67.010000 4.000000 ;
      END
   END in
   PIN out
      PORT
         LAYER met2 ;
	    RECT 46.110000 0.000000 46.740000 3.770000 ;
      END
   END out
   PIN pullupb
      PORT
         LAYER met2 ;
	    RECT 72.345000 0.000000 72.895000 3.770000 ;
      END
   END pullupb
   PIN pulldownb
      PORT
         LAYER met2 ;
	    RECT 62.750000 0.000000 63.305000 3.785000 ;
      END
   END pulldownb
   PIN outenb
      PORT
         LAYER met2 ;
	    RECT 50.345000 0.000000 50.900000 3.770000 ;
      END
   END outenb
   OBS
     LAYER li1 ;
       RECT 0.000000 4.000000 80.0000 165.0000 ;
     LAYER met1 ;
       RECT 0.000000 4.000000 80.0000 165.0000 ;
     LAYER met2 ;
       RECT 0.000000 4.000000 80.0000 165.0000 ;
     LAYER met3 ;
       RECT 0.000000 4.000000 80.0000 165.0000 ;
     LAYER met4 ;
       RECT 0.000000 4.000000 80.0000 165.0000 ;
     LAYER met5 ;
       RECT 0.000000 4.000000 80.0000 165.0000 ;
   END
END digital_out_pad
MACRO analog200ohm_pad
   CLASS BLOCK ;
   FOREIGN analog200ohm_pad ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 80.0000 BY 165.0000 ;
   OBS
     LAYER li1 ;
       RECT 0.000000 0.000000 80.0000 165.0000 ;
     LAYER met1 ;
       RECT 0.000000 0.000000 80.0000 165.0000 ;
     LAYER met2 ;
       RECT 0.000000 0.000000 80.0000 165.0000 ;
     LAYER met3 ;
       RECT 0.000000 0.000000 80.0000 165.0000 ;
     LAYER met4 ;
       RECT 0.000000 0.000000 80.0000 165.0000 ;
     LAYER met5 ;
       RECT 0.000000 0.000000 80.0000 165.0000 ;
   END
END analog200ohm_pad
MACRO vddio_pad
   CLASS BLOCK ;
   FOREIGN vddio_pad ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 80.0000 BY 165.0000 ;
   PIN VDD1V8
      PORT
         LAYER met5 ;
	    RECT 0.0000 0.0000 0.5000 5.0000 ;
      END
   END VDD1V8
   PIN VSS
      PORT
         LAYER met5 ;
	    RECT 0.0000 7.0000 0.5000 22.0000 ;
      END
   END VSS
   PIN VDD3V3
      PORT
         LAYER met5 ;
	    RECT 0.0000 24.0000 0.5000 39.0000 ;
      END
   END VDD3V3
   PIN VSSIO
      PORT
         LAYER met5 ;
	    RECT 0.0000 41.0000 0.5000 56.0000 ;
      END
   END VSSIO
   PIN VDDIO
      PORT
         LAYER met5 ;
	    RECT 12.9050 83.4650 66.4750 144.3350 ;
      END
   END VDDIO
   OBS
     LAYER li1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met2 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met3 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met4 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met5 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
   END
END vddio_pad
MACRO vdd1v8_pad
   CLASS BLOCK ;
   FOREIGN vdd1v8_pad ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 80.0000 BY 165.0000 ;
   PIN VDD1V8
      PORT
         LAYER met5 ;
	    RECT 0.0000 0.0000 0.5000 5.0000 ;
      END
   END VDD1V8
   PIN VSS
      PORT
         LAYER met5 ;
	    RECT 0.0000 7.0000 0.5000 22.0000 ;
      END
   END VSS
   PIN VDD3V3
      PORT
         LAYER met5 ;
	    RECT 0.0000 24.0000 0.5000 39.0000 ;
      END
   END VDD3V3
   PIN VSSIO
      PORT
         LAYER met5 ;
	    RECT 0.0000 41.0000 0.5000 56.0000 ;
      END
   END VSSIO
   PIN VDDIO
      PORT
         LAYER met5 ;
	    RECT 0.0000 58.0000 0.5000 73.0000 ;
      END
   END VDDIO
   OBS
     LAYER li1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met2 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met3 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met4 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met5 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
   END
END vdd1v8_pad
MACRO vss_pad
   CLASS BLOCK ;
   FOREIGN vss_pad ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 80.0000 BY 165.0000 ;
   PIN VDD1V8
      PORT
         LAYER met5 ;
	    RECT 0.0000 0.0000 0.5000 5.0000 ;
      END
   END VDD1V8
   PIN VSS
      PORT
         LAYER met5 ;
	    RECT 0.0000 7.0000 0.5000 22.0000 ;
      END
   END VSS
   PIN VDD3V3
      PORT
         LAYER met5 ;
	    RECT 0.0000 24.0000 0.5000 39.0000 ;
      END
   END VDD3V3
   PIN VSSIO
      PORT
         LAYER met5 ;
	    RECT 0.0000 41.0000 0.5000 56.0000 ;
      END
   END VSSIO
   PIN VDDIO
      PORT
         LAYER met5 ;
	    RECT 0.0000 58.0000 0.5000 73.0000 ;
      END
   END VDDIO
   OBS
     LAYER li1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met2 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met3 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met4 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met5 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
   END
END vss_pad
MACRO analog_pad
   CLASS BLOCK ;
   FOREIGN analog_pad ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 80.0000 BY 165.0000 ;
   OBS
     LAYER li1 ;
       RECT 0.000000 0.000000 80.0000 165.0000 ;
     LAYER met1 ;
       RECT 0.000000 0.000000 80.0000 165.0000 ;
     LAYER met2 ;
       RECT 0.000000 0.000000 80.0000 165.0000 ;
     LAYER met3 ;
       RECT 0.000000 0.000000 80.0000 165.0000 ;
     LAYER met4 ;
       RECT 0.000000 0.000000 80.0000 165.0000 ;
     LAYER met5 ;
       RECT 0.000000 0.000000 80.0000 165.0000 ;
   END
END analog_pad
MACRO pad_spacer_50um
   CLASS BLOCK ;
   FOREIGN pad_spacer_50um ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 50.0000 BY 165.0000 ;
   PIN VDD1V8
      PORT
         LAYER met5 ;
	    RECT 0.0000 0.0000 0.5000 5.0000 ;
      END
   END VDD1V8
   PIN VSS
      PORT
         LAYER met5 ;
	    RECT 0.0000 7.0000 0.5000 22.0000 ;
      END
   END VSS
   PIN VDD3V3
      PORT
         LAYER met5 ;
	    RECT 0.0000 24.0000 0.5000 39.0000 ;
      END
   END VDD3V3
   PIN VSSIO
      PORT
         LAYER met5 ;
	    RECT 0.0000 41.0000 0.5000 56.0000 ;
      END
   END VSSIO
   PIN VDDIO
      PORT
         LAYER met5 ;
	    RECT 0.0000 58.0000 0.5000 73.0000 ;
      END
   END VDDIO
   OBS
     LAYER li1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met2 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met3 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met4 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met5 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
   END
END pad_spacer_50um
MACRO pad_spacer_20um
   CLASS BLOCK ;
   FOREIGN pad_spacer_20um ;
   ORIGIN 0.0000 0.0000 ;
   SIZE 20.0000 BY 165.0000 ;
   OBS
   END
END pad_spacer_20um
MACRO pad_spacer_10um
   CLASS BLOCK ;
   FOREIGN pad_spacer_10um ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 10.0000 BY 165.0000 ;
   PIN VDD1V8
      PORT
         LAYER met5 ;
	    RECT 9.5000 0.0000 10.0000 5.0000 ;
      END
   END VDD1V8
   PIN VSS
      PORT
         LAYER met5 ;
	    RECT 9.5000 7.0000 10.0000 22.0000 ;
      END
   END VSS
   PIN VDD3V3
      PORT
         LAYER met5 ;
	    RECT 9.5000 24.0000 10.0000 39.0000 ;
      END
   END VDD3V3
   PIN VSSIO
      PORT
         LAYER met5 ;
	    RECT 9.3000 155.0000 10.0000 165.0000 ;
      END
   END VSSIO
   PIN VDDIO
      PORT
         LAYER met5 ;
	    RECT 9.5000 58.0000 10.0000 73.0000 ;
      END
   END VDDIO
   OBS
     LAYER li1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met2 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met3 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met4 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met5 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
   END
END pad_spacer_10um
MACRO pad_spacer_2um
   CLASS BLOCK ;
   FOREIGN pad_spacer_2um ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 2.0000 BY 165.0000 ;
   PIN VDD1V8
      PORT
         LAYER met5 ;
	    RECT 0.0000 0.0000 2.0000 5.0000 ;
      END
   END VDD1V8
   PIN VSS
      PORT
         LAYER met5 ;
	    RECT 0.0000 7.0000 2.0000 22.0000 ;
      END
   END VSS
   PIN VDD3V3
      PORT
         LAYER met5 ;
	    RECT 0.0000 24.0000 2.0000 39.0000 ;
      END
   END VDD3V3
   PIN VSSIO
      PORT
         LAYER met5 ;
	    RECT 0.0000 41.0000 2.0000 56.0000 ;
      END
   END VSSIO
   PIN VDDIO
      PORT
         LAYER met5 ;
	    RECT 0.0000 58.0000 2.0000 73.0000 ;
      END
   END VDDIO
   OBS
     LAYER li1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met2 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met3 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met4 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met5 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
   END
END pad_spacer_2um
MACRO pad_spacer_1um
   CLASS BLOCK ;
   FOREIGN pad_spacer_1um ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 1.0000 BY 165.0000 ;
   PIN VDD1V8
      PORT
         LAYER met5 ;
	    RECT -0.3000 0.0000 1.3000 5.0000 ;
      END
   END VDD1V8
   PIN VSS
      PORT
         LAYER met5 ;
	    RECT -0.3000 7.0000 1.3000 22.0000 ;
      END
   END VSS
   PIN VDD3V3
      PORT
         LAYER met5 ;
	    RECT -0.3000 24.0000 1.3000 39.0000 ;
      END
   END VDD3V3
   PIN VSSIO
      PORT
         LAYER met5 ;
	    RECT -0.3000 41.0000 1.3000 56.0000 ;
      END
   END VSSIO
   PIN VDDIO
      PORT
         LAYER met5 ;
	    RECT -0.3000 58.0000 1.3000 73.0000 ;
      END
   END VDDIO
   OBS
     LAYER li1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met2 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met3 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met4 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met5 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
   END
END pad_spacer_1um
MACRO vssio_pad
   CLASS BLOCK ;
   FOREIGN vssio_pad ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 80.0000 BY 165.0000 ;
   PIN VDD1V8
      PORT
         LAYER met5 ;
	    RECT 0.0000 0.0000 0.5000 5.0000 ;
      END
   END VDD1V8
   PIN VSS
      PORT
         LAYER met5 ;
	    RECT 0.0000 7.0000 0.5000 22.0000 ;
      END
   END VSS
   PIN VDD3V3
      PORT
         LAYER met5 ;
	    RECT 0.0000 24.0000 0.5000 39.0000 ;
      END
   END VDD3V3
   PIN VSSIO
      PORT
         LAYER met5 ;
	    RECT 0.0000 41.0000 0.5000 56.0000 ;
      END
   END VSSIO
   PIN VDDIO
      PORT
         LAYER met5 ;
	    RECT 0.0000 58.0000 0.5000 73.0000 ;
      END
   END VDDIO
   OBS
     LAYER li1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met2 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met3 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met4 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met5 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
   END
END vssio_pad
MACRO vdd3v3_pad
   CLASS BLOCK ;
   FOREIGN vdd3v3_pad ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 80.0000 BY 165.0000 ;
   PIN VDD1V8
      PORT
         LAYER met5 ;
	    RECT 0.0000 0.0000 0.5000 5.0000 ;
      END
   END VDD1V8
   PIN VSS
      PORT
         LAYER met5 ;
	    RECT 0.0000 7.0000 0.5000 22.0000 ;
      END
   END VSS
   PIN VDD3V3
      PORT
         LAYER met5 ;
	    RECT 0.0000 24.0000 0.5000 39.0000 ;
      END
   END VDD3V3
   PIN VSSIO
      PORT
         LAYER met5 ;
	    RECT 0.0000 41.0000 0.5000 56.0000 ;
      END
   END VSSIO
   PIN VDDIO
      PORT
         LAYER met5 ;
	    RECT 0.0000 58.0000 0.5000 73.0000 ;
      END
   END VDDIO
   OBS
     LAYER li1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met2 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met3 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met4 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met5 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
   END
END vdd3v3_pad
MACRO pad_spacer_5um
   CLASS BLOCK ;
   FOREIGN pad_spacer_5um ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.0000 BY 165.0000 ;
   PIN VDD1V8
      PORT
         LAYER met5 ;
	    RECT 4.5000 0.0000 5.0000 5.0000 ;
      END
   END VDD1V8
   PIN VSS
      PORT
         LAYER met5 ;
	    RECT 4.5000 7.0000 5.0000 22.0000 ;
      END
   END VSS
   PIN VDD3V3
      PORT
         LAYER met5 ;
	    RECT 4.5000 24.0000 5.0000 39.0000 ;
      END
   END VDD3V3
   PIN VSSIO
      PORT
         LAYER met5 ;
	    RECT 4.5000 41.0000 5.0000 56.0000 ;
      END
   END VSSIO
   PIN VDDIO
      PORT
         LAYER met5 ;
	    RECT 4.5000 58.0000 5.0000 73.0000 ;
      END
   END VDDIO
   OBS
     LAYER li1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met1 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met2 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met3 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met4 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
     LAYER met5 ;
       RECT 0.000000 0.000000 0.0 0.0 ;
   END
END pad_spacer_5um
MACRO digital_in_pad
   CLASS BLOCK ;
   FOREIGN digital_in_pad ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 80.0000 BY 165.0000 ;
   PIN in3v
      PORT
         LAYER met2 ;
	    RECT 63.890000 0.000000 64.930000 4.000000 ;
      END
   END in3v
   PIN in
      PORT
         LAYER met2 ;
	    RECT 65.920000 0.000000 66.960000 4.000000 ;
      END
   END in
   OBS
     LAYER li1 ;
       RECT 0.000000 4.000000 80.0000 165.0000 ;
     LAYER met1 ;
       RECT 0.000000 4.000000 80.0000 165.0000 ;
     LAYER met2 ;
       RECT 0.000000 4.000000 80.0000 165.0000 ;
     LAYER met3 ;
       RECT 0.000000 4.000000 80.0000 165.0000 ;
     LAYER met4 ;
       RECT 0.000000 4.000000 80.0000 165.0000 ;
     LAYER met5 ;
       RECT 0.000000 4.000000 80.0000 165.0000 ;
   END
END digital_in_pad
MACRO corner_pad
   CLASS BLOCK ;
   FOREIGN corner_pad ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 175.0000 BY 175.0000 ;
   OBS
     LAYER li1 ;
       RECT 0.000000 0.000000 175.0000 175.0000 ;
     LAYER met1 ;
       RECT 0.000000 0.000000 175.0000 175.0000 ;
     LAYER met2 ;
       RECT 0.000000 0.000000 175.0000 175.0000 ;
     LAYER met3 ;
       RECT 0.000000 0.000000 175.0000 175.0000 ;
     LAYER met4 ;
       RECT 0.000000 0.000000 175.0000 175.0000 ;
     LAYER met5 ;
       RECT 0.000000 0.000000 175.0000 175.0000 ;
   END
END corner_pad
END LIBRARY ;
