magic
tech sky130A
timestamp 1636140409
<< obsm1 >>
rect 62 62 68248 41592
<< obsm2 >>
rect 62 62 68248 41592
<< metal3 >>
rect 136 41344 68174 41518
rect 476 41004 67834 41178
rect 68204 39576 68310 39614
rect 0 18428 106 18466
rect 0 17952 106 17990
rect 0 16864 106 16902
rect 0 16388 106 16426
rect 0 15504 106 15542
rect 0 14960 106 14998
rect 0 14076 106 14114
rect 68204 9656 68310 9694
rect 68204 8840 68310 8878
rect 68204 8160 68310 8198
rect 68204 7412 68310 7450
rect 68204 6800 68310 6838
rect 0 4964 106 5002
rect 0 4148 106 4186
rect 0 4012 106 4050
rect 476 476 67834 650
rect 136 136 68174 310
<< obsm3 >>
rect 62 41578 68248 41592
rect 62 41284 76 41578
rect 68234 41284 68248 41578
rect 62 41238 68248 41284
rect 62 40944 416 41238
rect 67894 40944 68248 41238
rect 62 39674 68248 40944
rect 62 39516 68144 39674
rect 62 18526 68248 39516
rect 166 18368 68248 18526
rect 62 18050 68248 18368
rect 166 17892 68248 18050
rect 62 16962 68248 17892
rect 166 16804 68248 16962
rect 62 16486 68248 16804
rect 166 16328 68248 16486
rect 62 15602 68248 16328
rect 166 15444 68248 15602
rect 62 15058 68248 15444
rect 166 14900 68248 15058
rect 62 14174 68248 14900
rect 166 14016 68248 14174
rect 62 9754 68248 14016
rect 62 9596 68144 9754
rect 62 8938 68248 9596
rect 62 8780 68144 8938
rect 62 8258 68248 8780
rect 62 8100 68144 8258
rect 62 7510 68248 8100
rect 62 7352 68144 7510
rect 62 6898 68248 7352
rect 62 6740 68144 6898
rect 62 5062 68248 6740
rect 166 4904 68248 5062
rect 62 4246 68248 4904
rect 166 3952 68248 4246
rect 62 710 68248 3952
rect 62 416 416 710
rect 67894 416 68248 710
rect 62 370 68248 416
rect 62 76 76 370
rect 68234 76 68248 370
rect 62 62 68248 76
<< metal4 >>
rect 136 136 310 41518
rect 14348 41548 14386 41654
rect 15504 41548 15542 41654
rect 16728 41548 16766 41654
rect 18088 41548 18126 41654
rect 19244 41548 19282 41654
rect 20536 41548 20574 41654
rect 21760 41548 21798 41654
rect 23052 41548 23090 41654
rect 24276 41548 24314 41654
rect 25568 41548 25606 41654
rect 26792 41548 26830 41654
rect 28084 41548 28122 41654
rect 29240 41548 29278 41654
rect 30464 41548 30502 41654
rect 31824 41548 31862 41654
rect 33048 41548 33086 41654
rect 34272 41548 34310 41654
rect 35496 41548 35534 41654
rect 36788 41548 36826 41654
rect 37944 41548 37982 41654
rect 39304 41548 39342 41654
rect 40528 41548 40566 41654
rect 41752 41548 41790 41654
rect 42976 41548 43014 41654
rect 44200 41548 44238 41654
rect 45492 41548 45530 41654
rect 46784 41548 46822 41654
rect 48008 41548 48046 41654
rect 49232 41548 49270 41654
rect 50524 41548 50562 41654
rect 51680 41548 51718 41654
rect 53040 41548 53078 41654
rect 59228 41548 59266 41654
rect 59840 41548 59878 41654
rect 65416 41548 65454 41654
rect 476 476 650 41178
rect 67660 476 67834 41178
rect 8024 0 8062 106
rect 8568 0 8606 106
rect 9112 0 9150 106
rect 9792 0 9830 106
rect 10268 0 10306 106
rect 10880 0 10918 106
rect 11560 0 11598 106
rect 12104 0 12142 106
rect 12716 0 12754 106
rect 13260 0 13298 106
rect 13804 0 13842 106
rect 14144 0 14182 106
rect 14348 0 14386 106
rect 15028 0 15066 106
rect 15368 0 15406 106
rect 15640 0 15678 106
rect 16184 0 16222 106
rect 16728 0 16766 106
rect 16796 0 16834 106
rect 17272 0 17310 106
rect 17952 0 17990 106
rect 18020 0 18058 106
rect 18496 0 18534 106
rect 19040 0 19078 106
rect 19244 0 19282 106
rect 19720 0 19758 106
rect 20332 0 20370 106
rect 20536 0 20574 106
rect 20876 0 20914 106
rect 21420 0 21458 106
rect 21760 0 21798 106
rect 21964 0 22002 106
rect 22644 0 22682 106
rect 22984 0 23022 106
rect 23188 0 23226 106
rect 23800 0 23838 106
rect 24140 0 24178 106
rect 24344 0 24382 106
rect 24888 0 24926 106
rect 25500 0 25538 106
rect 25568 0 25606 106
rect 26112 0 26150 106
rect 26656 0 26694 106
rect 26792 0 26830 106
rect 27200 0 27238 106
rect 27880 0 27918 106
rect 28016 0 28054 106
rect 28492 0 28530 106
rect 29036 0 29074 106
rect 29240 0 29278 106
rect 29580 0 29618 106
rect 30464 0 30502 106
rect 31756 0 31794 106
rect 32980 0 33018 106
rect 34136 0 34174 106
rect 35496 0 35534 106
rect 36720 0 36758 106
rect 37944 0 37982 106
rect 39236 0 39274 106
rect 40460 0 40498 106
rect 41752 0 41790 106
rect 42976 0 43014 106
rect 44268 0 44306 106
rect 45492 0 45530 106
rect 46716 0 46754 106
rect 47940 0 47978 106
rect 49232 0 49270 106
rect 50456 0 50494 106
rect 51680 0 51718 106
rect 52972 0 53010 106
rect 61608 0 61646 106
rect 61676 0 61714 106
rect 68000 136 68174 41518
<< obsm4 >>
rect 62 41578 14288 41592
rect 62 76 76 41578
rect 370 41488 14288 41578
rect 14446 41488 15444 41592
rect 15602 41488 16668 41592
rect 16826 41488 18028 41592
rect 18186 41488 19184 41592
rect 19342 41488 20476 41592
rect 20634 41488 21700 41592
rect 21858 41488 22992 41592
rect 23150 41488 24216 41592
rect 24374 41488 25508 41592
rect 25666 41488 26732 41592
rect 26890 41488 28024 41592
rect 28182 41488 29180 41592
rect 29338 41488 30404 41592
rect 30562 41488 31764 41592
rect 31922 41488 32988 41592
rect 33146 41488 34212 41592
rect 34370 41488 35436 41592
rect 35594 41488 36728 41592
rect 36886 41488 37884 41592
rect 38042 41488 39244 41592
rect 39402 41488 40468 41592
rect 40626 41488 41692 41592
rect 41850 41488 42916 41592
rect 43074 41488 44140 41592
rect 44298 41488 45432 41592
rect 45590 41488 46724 41592
rect 46882 41488 47948 41592
rect 48106 41488 49172 41592
rect 49330 41488 50464 41592
rect 50622 41488 51620 41592
rect 51778 41488 52980 41592
rect 53138 41488 59168 41592
rect 59326 41488 59780 41592
rect 59938 41488 65356 41592
rect 65514 41578 68248 41592
rect 65514 41488 67940 41578
rect 370 41238 67940 41488
rect 370 416 416 41238
rect 710 416 67600 41238
rect 67894 416 67940 41238
rect 370 166 67940 416
rect 370 76 7964 166
rect 62 62 7964 76
rect 8122 62 8508 166
rect 8666 62 9052 166
rect 9210 62 9732 166
rect 9890 62 10208 166
rect 10366 62 10820 166
rect 10978 62 11500 166
rect 11658 62 12044 166
rect 12202 62 12656 166
rect 12814 62 13200 166
rect 13358 62 13744 166
rect 13902 62 14084 166
rect 14242 62 14288 166
rect 14446 62 14968 166
rect 15126 62 15308 166
rect 15466 62 15580 166
rect 15738 62 16124 166
rect 16282 62 16668 166
rect 16894 62 17212 166
rect 17370 62 17892 166
rect 18118 62 18436 166
rect 18594 62 18980 166
rect 19138 62 19184 166
rect 19342 62 19660 166
rect 19818 62 20272 166
rect 20430 62 20476 166
rect 20634 62 20816 166
rect 20974 62 21360 166
rect 21518 62 21700 166
rect 21858 62 21904 166
rect 22062 62 22584 166
rect 22742 62 22924 166
rect 23082 62 23128 166
rect 23286 62 23740 166
rect 23898 62 24080 166
rect 24238 62 24284 166
rect 24442 62 24828 166
rect 24986 62 25440 166
rect 25666 62 26052 166
rect 26210 62 26596 166
rect 26890 62 27140 166
rect 27298 62 27820 166
rect 28114 62 28432 166
rect 28590 62 28976 166
rect 29134 62 29180 166
rect 29338 62 29520 166
rect 29678 62 30404 166
rect 30562 62 31696 166
rect 31854 62 32920 166
rect 33078 62 34076 166
rect 34234 62 35436 166
rect 35594 62 36660 166
rect 36818 62 37884 166
rect 38042 62 39176 166
rect 39334 62 40400 166
rect 40558 62 41692 166
rect 41850 62 42916 166
rect 43074 62 44208 166
rect 44366 62 45432 166
rect 45590 62 46656 166
rect 46814 62 47880 166
rect 48038 62 49172 166
rect 49330 62 50396 166
rect 50554 62 51620 166
rect 51778 62 52912 166
rect 53070 62 61548 166
rect 61774 76 67940 166
rect 68234 76 68248 41578
rect 61774 62 68248 76
<< labels >>
rlabel metal4 s 11560 0 11598 106 6 din0[0]
port 1 nsew default input
rlabel metal4 s 12104 0 12142 106 6 din0[1]
port 2 nsew default input
rlabel metal4 s 12716 0 12754 106 6 din0[2]
port 3 nsew default input
rlabel metal4 s 13260 0 13298 106 6 din0[3]
port 4 nsew default input
rlabel metal4 s 13804 0 13842 106 6 din0[4]
port 5 nsew default input
rlabel metal4 s 14348 0 14386 106 6 din0[5]
port 6 nsew default input
rlabel metal4 s 15028 0 15066 106 6 din0[6]
port 7 nsew default input
rlabel metal4 s 15640 0 15678 106 6 din0[7]
port 8 nsew default input
rlabel metal4 s 16184 0 16222 106 6 din0[8]
port 9 nsew default input
rlabel metal4 s 16728 0 16766 106 6 din0[9]
port 10 nsew default input
rlabel metal4 s 17272 0 17310 106 6 din0[10]
port 11 nsew default input
rlabel metal4 s 17952 0 17990 106 6 din0[11]
port 12 nsew default input
rlabel metal4 s 18496 0 18534 106 6 din0[12]
port 13 nsew default input
rlabel metal4 s 19040 0 19078 106 6 din0[13]
port 14 nsew default input
rlabel metal4 s 19720 0 19758 106 6 din0[14]
port 15 nsew default input
rlabel metal4 s 20332 0 20370 106 6 din0[15]
port 16 nsew default input
rlabel metal4 s 20876 0 20914 106 6 din0[16]
port 17 nsew default input
rlabel metal4 s 21420 0 21458 106 6 din0[17]
port 18 nsew default input
rlabel metal4 s 21964 0 22002 106 6 din0[18]
port 19 nsew default input
rlabel metal4 s 22644 0 22682 106 6 din0[19]
port 20 nsew default input
rlabel metal4 s 23188 0 23226 106 6 din0[20]
port 21 nsew default input
rlabel metal4 s 23800 0 23838 106 6 din0[21]
port 22 nsew default input
rlabel metal4 s 24344 0 24382 106 6 din0[22]
port 23 nsew default input
rlabel metal4 s 24888 0 24926 106 6 din0[23]
port 24 nsew default input
rlabel metal4 s 25568 0 25606 106 6 din0[24]
port 25 nsew default input
rlabel metal4 s 26112 0 26150 106 6 din0[25]
port 26 nsew default input
rlabel metal4 s 26656 0 26694 106 6 din0[26]
port 27 nsew default input
rlabel metal4 s 27200 0 27238 106 6 din0[27]
port 28 nsew default input
rlabel metal4 s 27880 0 27918 106 6 din0[28]
port 29 nsew default input
rlabel metal4 s 28492 0 28530 106 6 din0[29]
port 30 nsew default input
rlabel metal4 s 29036 0 29074 106 6 din0[30]
port 31 nsew default input
rlabel metal4 s 29580 0 29618 106 6 din0[31]
port 32 nsew default input
rlabel metal4 s 8024 0 8062 106 6 addr0[0]
port 33 nsew default input
rlabel metal4 s 8568 0 8606 106 6 addr0[1]
port 34 nsew default input
rlabel metal3 s 0 14076 106 14114 6 addr0[2]
port 35 nsew default input
rlabel metal3 s 0 14960 106 14998 6 addr0[3]
port 36 nsew default input
rlabel metal3 s 0 15504 106 15542 6 addr0[4]
port 37 nsew default input
rlabel metal3 s 0 16388 106 16426 6 addr0[5]
port 38 nsew default input
rlabel metal3 s 0 16864 106 16902 6 addr0[6]
port 39 nsew default input
rlabel metal3 s 0 17952 106 17990 6 addr0[7]
port 40 nsew default input
rlabel metal3 s 0 18428 106 18466 6 addr0[8]
port 41 nsew default input
rlabel metal4 s 59840 41548 59878 41654 6 addr1[0]
port 42 nsew default input
rlabel metal4 s 59228 41548 59266 41654 6 addr1[1]
port 43 nsew default input
rlabel metal3 s 68204 9656 68310 9694 6 addr1[2]
port 44 nsew default input
rlabel metal3 s 68204 8840 68310 8878 6 addr1[3]
port 45 nsew default input
rlabel metal3 s 68204 8160 68310 8198 6 addr1[4]
port 46 nsew default input
rlabel metal3 s 68204 7412 68310 7450 6 addr1[5]
port 47 nsew default input
rlabel metal3 s 68204 6800 68310 6838 6 addr1[6]
port 48 nsew default input
rlabel metal4 s 61608 0 61646 106 6 addr1[7]
port 49 nsew default input
rlabel metal4 s 61676 0 61714 106 6 addr1[8]
port 50 nsew default input
rlabel metal3 s 0 4012 106 4050 6 csb0
port 51 nsew default input
rlabel metal3 s 68204 39576 68310 39614 6 csb1
port 52 nsew default input
rlabel metal3 s 0 4964 106 5002 6 web0
port 53 nsew default input
rlabel metal3 s 0 4148 106 4186 6 clk0
port 54 nsew default input
rlabel metal4 s 65416 41548 65454 41654 6 clk1
port 55 nsew default input
rlabel metal4 s 9112 0 9150 106 6 wmask0[0]
port 56 nsew default input
rlabel metal4 s 9792 0 9830 106 6 wmask0[1]
port 57 nsew default input
rlabel metal4 s 10268 0 10306 106 6 wmask0[2]
port 58 nsew default input
rlabel metal4 s 10880 0 10918 106 6 wmask0[3]
port 59 nsew default input
rlabel metal4 s 14144 0 14182 106 6 dout0[0]
port 60 nsew default output
rlabel metal4 s 15368 0 15406 106 6 dout0[1]
port 61 nsew default output
rlabel metal4 s 16796 0 16834 106 6 dout0[2]
port 62 nsew default output
rlabel metal4 s 18020 0 18058 106 6 dout0[3]
port 63 nsew default output
rlabel metal4 s 19244 0 19282 106 6 dout0[4]
port 64 nsew default output
rlabel metal4 s 20536 0 20574 106 6 dout0[5]
port 65 nsew default output
rlabel metal4 s 21760 0 21798 106 6 dout0[6]
port 66 nsew default output
rlabel metal4 s 22984 0 23022 106 6 dout0[7]
port 67 nsew default output
rlabel metal4 s 24140 0 24178 106 6 dout0[8]
port 68 nsew default output
rlabel metal4 s 25500 0 25538 106 6 dout0[9]
port 69 nsew default output
rlabel metal4 s 26792 0 26830 106 6 dout0[10]
port 70 nsew default output
rlabel metal4 s 28016 0 28054 106 6 dout0[11]
port 71 nsew default output
rlabel metal4 s 29240 0 29278 106 6 dout0[12]
port 72 nsew default output
rlabel metal4 s 30464 0 30502 106 6 dout0[13]
port 73 nsew default output
rlabel metal4 s 31756 0 31794 106 6 dout0[14]
port 74 nsew default output
rlabel metal4 s 32980 0 33018 106 6 dout0[15]
port 75 nsew default output
rlabel metal4 s 34136 0 34174 106 6 dout0[16]
port 76 nsew default output
rlabel metal4 s 35496 0 35534 106 6 dout0[17]
port 77 nsew default output
rlabel metal4 s 36720 0 36758 106 6 dout0[18]
port 78 nsew default output
rlabel metal4 s 37944 0 37982 106 6 dout0[19]
port 79 nsew default output
rlabel metal4 s 39236 0 39274 106 6 dout0[20]
port 80 nsew default output
rlabel metal4 s 40460 0 40498 106 6 dout0[21]
port 81 nsew default output
rlabel metal4 s 41752 0 41790 106 6 dout0[22]
port 82 nsew default output
rlabel metal4 s 42976 0 43014 106 6 dout0[23]
port 83 nsew default output
rlabel metal4 s 44268 0 44306 106 6 dout0[24]
port 84 nsew default output
rlabel metal4 s 45492 0 45530 106 6 dout0[25]
port 85 nsew default output
rlabel metal4 s 46716 0 46754 106 6 dout0[26]
port 86 nsew default output
rlabel metal4 s 47940 0 47978 106 6 dout0[27]
port 87 nsew default output
rlabel metal4 s 49232 0 49270 106 6 dout0[28]
port 88 nsew default output
rlabel metal4 s 50456 0 50494 106 6 dout0[29]
port 89 nsew default output
rlabel metal4 s 51680 0 51718 106 6 dout0[30]
port 90 nsew default output
rlabel metal4 s 52972 0 53010 106 6 dout0[31]
port 91 nsew default output
rlabel metal4 s 14348 41548 14386 41654 6 dout1[0]
port 92 nsew default output
rlabel metal4 s 15504 41548 15542 41654 6 dout1[1]
port 93 nsew default output
rlabel metal4 s 16728 41548 16766 41654 6 dout1[2]
port 94 nsew default output
rlabel metal4 s 18088 41548 18126 41654 6 dout1[3]
port 95 nsew default output
rlabel metal4 s 19244 41548 19282 41654 6 dout1[4]
port 96 nsew default output
rlabel metal4 s 20536 41548 20574 41654 6 dout1[5]
port 97 nsew default output
rlabel metal4 s 21760 41548 21798 41654 6 dout1[6]
port 98 nsew default output
rlabel metal4 s 23052 41548 23090 41654 6 dout1[7]
port 99 nsew default output
rlabel metal4 s 24276 41548 24314 41654 6 dout1[8]
port 100 nsew default output
rlabel metal4 s 25568 41548 25606 41654 6 dout1[9]
port 101 nsew default output
rlabel metal4 s 26792 41548 26830 41654 6 dout1[10]
port 102 nsew default output
rlabel metal4 s 28084 41548 28122 41654 6 dout1[11]
port 103 nsew default output
rlabel metal4 s 29240 41548 29278 41654 6 dout1[12]
port 104 nsew default output
rlabel metal4 s 30464 41548 30502 41654 6 dout1[13]
port 105 nsew default output
rlabel metal4 s 31824 41548 31862 41654 6 dout1[14]
port 106 nsew default output
rlabel metal4 s 33048 41548 33086 41654 6 dout1[15]
port 107 nsew default output
rlabel metal4 s 34272 41548 34310 41654 6 dout1[16]
port 108 nsew default output
rlabel metal4 s 35496 41548 35534 41654 6 dout1[17]
port 109 nsew default output
rlabel metal4 s 36788 41548 36826 41654 6 dout1[18]
port 110 nsew default output
rlabel metal4 s 37944 41548 37982 41654 6 dout1[19]
port 111 nsew default output
rlabel metal4 s 39304 41548 39342 41654 6 dout1[20]
port 112 nsew default output
rlabel metal4 s 40528 41548 40566 41654 6 dout1[21]
port 113 nsew default output
rlabel metal4 s 41752 41548 41790 41654 6 dout1[22]
port 114 nsew default output
rlabel metal4 s 42976 41548 43014 41654 6 dout1[23]
port 115 nsew default output
rlabel metal4 s 44200 41548 44238 41654 6 dout1[24]
port 116 nsew default output
rlabel metal4 s 45492 41548 45530 41654 6 dout1[25]
port 117 nsew default output
rlabel metal4 s 46784 41548 46822 41654 6 dout1[26]
port 118 nsew default output
rlabel metal4 s 48008 41548 48046 41654 6 dout1[27]
port 119 nsew default output
rlabel metal4 s 49232 41548 49270 41654 6 dout1[28]
port 120 nsew default output
rlabel metal4 s 50524 41548 50562 41654 6 dout1[29]
port 121 nsew default output
rlabel metal4 s 51680 41548 51718 41654 6 dout1[30]
port 122 nsew default output
rlabel metal4 s 53040 41548 53078 41654 6 dout1[31]
port 123 nsew default output
rlabel metal3 s 476 476 67834 650 6 vccd1
port 124 nsew power bidirectional abutment
rlabel metal3 s 476 41004 67834 41178 6 vccd1
port 124 nsew power bidirectional abutment
rlabel metal4 s 67660 476 67834 41178 6 vccd1
port 124 nsew power bidirectional abutment
rlabel metal4 s 476 476 650 41178 6 vccd1
port 124 nsew power bidirectional abutment
rlabel metal3 s 136 41344 68174 41518 6 vssd1
port 125 nsew ground bidirectional abutment
rlabel metal3 s 136 136 68174 310 6 vssd1
port 125 nsew ground bidirectional abutment
rlabel metal4 s 136 136 310 41518 6 vssd1
port 125 nsew ground bidirectional abutment
rlabel metal4 s 68000 136 68174 41518 6 vssd1
port 125 nsew ground bidirectional abutment
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 68310 41654
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_END 15213044
string GDS_START 13196574
<< end >>
