VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS
MACRO digital_pll
   CLASS BLOCK ;
   FOREIGN digital_pll ;
   ORIGIN 0.000000 0.000000 ;
   SIZE 122.0300 BY 122.0300 ;
   PIN reset
      DIRECTION INPUT ;
      PORT
         LAYER met2 ;
	    RECT 72.950000 117.910000 73.510000 122.030000 ;
      END
   END reset
   PIN osc
      DIRECTION INPUT ;
      PORT
         LAYER met2 ;
	    RECT 3.950000 0.000000 4.510000 4.120000 ;
      END
   END osc
   PIN clockp[1]
      DIRECTION OUTPUT TRISTATE ;
      PORT
         LAYER met3 ;
	    RECT 0.000000 89.420000 4.200000 90.620000 ;
      END
   END clockp[1]
   PIN clockp[0]
      DIRECTION OUTPUT TRISTATE ;
      PORT
         LAYER met2 ;
	    RECT 43.510000 117.910000 44.070000 122.030000 ;
      END
   END clockp[0]
   PIN clockd[3]
      DIRECTION OUTPUT TRISTATE ;
      PORT
         LAYER met3 ;
	    RECT 0.000000 45.900000 4.200000 47.100000 ;
      END
   END clockd[3]
   PIN clockd[2]
      DIRECTION OUTPUT TRISTATE ;
      PORT
         LAYER met2 ;
	    RECT 62.830000 0.000000 63.390000 4.120000 ;
      END
   END clockd[2]
   PIN clockd[1]
      DIRECTION OUTPUT TRISTATE ;
      PORT
         LAYER met2 ;
	    RECT 92.270000 0.000000 92.830000 4.120000 ;
      END
   END clockd[1]
   PIN clockd[0]
      DIRECTION OUTPUT TRISTATE ;
      PORT
         LAYER met3 ;
	    RECT 117.830000 96.220000 122.030000 97.420000 ;
      END
   END clockd[0]
   PIN div[4]
      DIRECTION INPUT ;
      PORT
         LAYER met2 ;
	    RECT 14.070000 117.910000 14.630000 122.030000 ;
      END
   END div[4]
   PIN div[3]
      DIRECTION INPUT ;
      PORT
         LAYER met2 ;
	    RECT 33.390000 0.000000 33.950000 4.120000 ;
      END
   END div[3]
   PIN div[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
	    RECT 117.830000 9.180000 122.030000 10.380000 ;
      END
   END div[2]
   PIN div[1]
      DIRECTION INPUT ;
      PORT
         LAYER met2 ;
	    RECT 102.390000 117.910000 102.950000 122.030000 ;
      END
   END div[1]
   PIN div[0]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
	    RECT 117.830000 52.700000 122.030000 53.900000 ;
      END
   END div[0]
   OBS
         LAYER li1 ;
	    RECT 0.000000 0.000000 0 0 ;
   END
END digital_pll
