magic
tech sky130A
magscale 1 2
timestamp 1636140361
<< checkpaint >>
rect -1296 -1277 1772 2731
<< nwell >>
rect -36 679 512 1471
<< pwell >>
rect 340 25 442 159
<< psubdiff >>
rect 366 109 416 133
rect 366 75 374 109
rect 408 75 416 109
rect 366 51 416 75
<< nsubdiff >>
rect 366 1339 416 1363
rect 366 1305 374 1339
rect 408 1305 416 1339
rect 366 1281 416 1305
<< psubdiffcont >>
rect 374 75 408 109
<< nsubdiffcont >>
rect 374 1305 408 1339
<< poly >>
rect 114 703 144 907
rect 48 687 144 703
rect 48 653 64 687
rect 98 653 144 687
rect 48 637 144 653
rect 114 359 144 637
<< polycont >>
rect 64 653 98 687
<< locali >>
rect 0 1397 476 1431
rect 62 1130 96 1397
rect 64 687 98 703
rect 64 637 98 653
rect 166 687 200 1196
rect 270 1130 304 1397
rect 374 1339 408 1397
rect 374 1289 408 1305
rect 166 653 217 687
rect 166 144 200 653
rect 62 17 96 144
rect 270 17 304 144
rect 374 109 408 125
rect 374 17 408 75
rect 0 -17 476 17
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_16  sky130_sram_2kbyte_1rw1r_32x512_8_contact_16_0
timestamp 1636140361
transform 1 0 48 0 1 637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_29  sky130_sram_2kbyte_1rw1r_32x512_8_contact_29_0
timestamp 1636140361
transform 1 0 366 0 1 51
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_28  sky130_sram_2kbyte_1rw1r_32x512_8_contact_28_0
timestamp 1636140361
transform 1 0 366 0 1 1281
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m2_w1_260_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m2_w1_260_sli_dli_da_p_0
timestamp 1636140361
transform 1 0 54 0 1 51
box -26 -26 284 308
use sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m2_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m2_w2_000_sli_dli_da_p_0
timestamp 1636140361
transform 1 0 54 0 1 963
box -59 -56 317 454
<< labels >>
rlabel locali s 81 670 81 670 4 A
port 1 nsew
rlabel locali s 200 670 200 670 4 Z
port 2 nsew
rlabel locali s 238 0 238 0 4 gnd
port 3 nsew
rlabel locali s 238 1414 238 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 476 1414
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_END 392406
string GDS_START 390408
<< end >>
