module prim_lfsr (
	clk_i,
	rst_ni,
	seed_en_i,
	seed_i,
	lfsr_en_i,
	entropy_i,
	state_o
);
	parameter _sv2v_width_LfsrType = 56;
	parameter [_sv2v_width_LfsrType - 1:0] LfsrType = "GAL_XOR";
	parameter [31:0] LfsrDw = 32;
	parameter [31:0] EntropyDw = 8;
	parameter [31:0] StateOutDw = 8;
	function automatic signed [LfsrDw - 1:0] sv2v_cast_FFBD2_signed;
		input reg signed [LfsrDw - 1:0] inp;
		sv2v_cast_FFBD2_signed = inp;
	endfunction
	parameter [LfsrDw - 1:0] DefaultSeed = sv2v_cast_FFBD2_signed(1);
	parameter [LfsrDw - 1:0] CustomCoeffs = 1'sb0;
	parameter [0:0] MaxLenSVA = 1'b1;
	parameter [0:0] LockupSVA = 1'b1;
	parameter [0:0] ExtSeedSVA = 1'b1;
	input clk_i;
	input rst_ni;
	input seed_en_i;
	input [LfsrDw - 1:0] seed_i;
	input lfsr_en_i;
	input [EntropyDw - 1:0] entropy_i;
	output wire [StateOutDw - 1:0] state_o;
	localparam [31:0] GAL_XOR_LUT_OFF = 4;
	localparam [3903:0] GAL_XOR_COEFFS = {64'h0000000000000009, 64'h0000000000000012, 64'h0000000000000021, 64'h0000000000000041, 64'h000000000000008e, 64'h0000000000000108, 64'h0000000000000204, 64'h0000000000000402, 64'h0000000000000829, 64'h000000000000100d, 64'h0000000000002015, 64'h0000000000004001, 64'h0000000000008016, 64'h0000000000010004, 64'h0000000000020013, 64'h0000000000040013, 64'h0000000000080004, 64'h0000000000100002, 64'h0000000000200001, 64'h0000000000400010, 64'h000000000080000d, 64'h0000000001000004, 64'h0000000002000023, 64'h0000000004000013, 64'h0000000008000004, 64'h0000000010000002, 64'h0000000020000029, 64'h0000000040000004, 64'h0000000080000057, 64'h0000000100000029, 64'h0000000200000073, 64'h0000000400000002, 64'h000000080000003b, 64'h000000100000001f, 64'h0000002000000031, 64'h0000004000000008, 64'h000000800000001c, 64'h0000010000000004, 64'h000002000000001f, 64'h000004000000002c, 64'h0000080000000032, 64'h000010000000000d, 64'h0000200000000097, 64'h0000400000000010, 64'h000080000000005b, 64'h0001000000000038, 64'h000200000000000e, 64'h0004000000000025, 64'h0008000000000004, 64'h0010000000000023, 64'h002000000000003e, 64'h0040000000000023, 64'h008000000000004a, 64'h0100000000000016, 64'h0200000000000031, 64'h040000000000003d, 64'h0800000000000001, 64'h1000000000000013, 64'h2000000000000034, 64'h4000000000000001, 64'h800000000000000d};
	localparam [31:0] FIB_XNOR_LUT_OFF = 3;
	localparam [27887:0] FIB_XNOR_COEFFS = {168'h000000000000000000000000000000000000000006, 168'h00000000000000000000000000000000000000000c, 168'h000000000000000000000000000000000000000014, 168'h000000000000000000000000000000000000000030, 168'h000000000000000000000000000000000000000060, 168'h0000000000000000000000000000000000000000b8, 168'h000000000000000000000000000000000000000110, 168'h000000000000000000000000000000000000000240, 168'h000000000000000000000000000000000000000500, 168'h000000000000000000000000000000000000000829, 168'h00000000000000000000000000000000000000100d, 168'h000000000000000000000000000000000000002015, 168'h000000000000000000000000000000000000006000, 168'h00000000000000000000000000000000000000d008, 168'h000000000000000000000000000000000000012000, 168'h000000000000000000000000000000000000020400, 168'h000000000000000000000000000000000000040023, 168'h000000000000000000000000000000000000090000, 168'h000000000000000000000000000000000000140000, 168'h000000000000000000000000000000000000300000, 168'h000000000000000000000000000000000000420000, 168'h000000000000000000000000000000000000e10000, 168'h000000000000000000000000000000000001200000, 168'h000000000000000000000000000000000002000023, 168'h000000000000000000000000000000000004000013, 168'h000000000000000000000000000000000009000000, 168'h000000000000000000000000000000000014000000, 168'h000000000000000000000000000000000020000029, 168'h000000000000000000000000000000000048000000, 168'h000000000000000000000000000000000080200003, 168'h000000000000000000000000000000000100080000, 168'h000000000000000000000000000000000204000003, 168'h000000000000000000000000000000000500000000, 168'h000000000000000000000000000000000801000000, 168'h00000000000000000000000000000000100000001f, 168'h000000000000000000000000000000002000000031, 168'h000000000000000000000000000000004400000000, 168'h00000000000000000000000000000000a000140000, 168'h000000000000000000000000000000012000000000, 168'h0000000000000000000000000000000300000c0000, 168'h000000000000000000000000000000063000000000, 168'h0000000000000000000000000000000c0000030000, 168'h0000000000000000000000000000001b0000000000, 168'h000000000000000000000000000000300003000000, 168'h000000000000000000000000000000420000000000, 168'h000000000000000000000000000000c00000180000, 168'h000000000000000000000000000001008000000000, 168'h000000000000000000000000000003000000c00000, 168'h000000000000000000000000000006000c00000000, 168'h000000000000000000000000000009000000000000, 168'h000000000000000000000000000018003000000000, 168'h000000000000000000000000000030000000030000, 168'h000000000000000000000000000040000040000000, 168'h0000000000000000000000000000c0000600000000, 168'h000000000000000000000000000102000000000000, 168'h000000000000000000000000000200004000000000, 168'h000000000000000000000000000600003000000000, 168'h000000000000000000000000000c00000000000000, 168'h000000000000000000000000001800300000000000, 168'h000000000000000000000000003000000000000030, 168'h000000000000000000000000006000000000000000, 168'h00000000000000000000000000d800000000000000, 168'h000000000000000000000000010000400000000000, 168'h000000000000000000000000030180000000000000, 168'h000000000000000000000000060300000000000000, 168'h000000000000000000000000080400000000000000, 168'h000000000000000000000000140000028000000000, 168'h000000000000000000000000300060000000000000, 168'h000000000000000000000000410000000000000000, 168'h000000000000000000000000820000000001040000, 168'h000000000000000000000001000000800000000000, 168'h000000000000000000000003000600000000000000, 168'h000000000000000000000006018000000000000000, 168'h00000000000000000000000c000000018000000000, 168'h000000000000000000000018000000600000000000, 168'h000000000000000000000030000600000000000000, 168'h000000000000000000000040200000000000000000, 168'h0000000000000000000000c0000000060000000000, 168'h000000000000000000000110000000000000000000, 168'h000000000000000000000240000000480000000000, 168'h000000000000000000000600000000003000000000, 168'h000000000000000000000800400000000000000000, 168'h000000000000000000001800000300000000000000, 168'h000000000000000000003003000000000000000000, 168'h000000000000000000004002000000000000000000, 168'h00000000000000000000c000000000000000018000, 168'h000000000000000000010000000004000000000000, 168'h000000000000000000030000c00000000000000000, 168'h0000000000000000000600000000000000000000c0, 168'h0000000000000000000c00c0000000000000000000, 168'h000000000000000000140000000000000000000000, 168'h000000000000000000200001000000000000000000, 168'h000000000000000000400800000000000000000000, 168'h000000000000000000a00000000001400000000000, 168'h000000000000000001040000000000000000000000, 168'h000000000000000002004000000000000000000000, 168'h000000000000000005000000000028000000000000, 168'h000000000000000008000000004000000000000000, 168'h000000000000000018600000000000000000000000, 168'h000000000000000030000000000000000c00000000, 168'h000000000000000040200000000000000000000000, 168'h0000000000000000c0300000000000000000000000, 168'h000000000000000100010000000000000000000000, 168'h000000000000000200040000000000000000000000, 168'h0000000000000005000000000000000a0000000000, 168'h000000000000000800000010000000000000000000, 168'h000000000000001860000000000000000000000000, 168'h000000000000003003000000000000000000000000, 168'h000000000000004010000000000000000000000000, 168'h00000000000000a000000000140000000000000000, 168'h000000000000010080000000000000000000000000, 168'h000000000000030000000000000000000180000000, 168'h000000000000060018000000000000000000000000, 168'h0000000000000c0000000000000000300000000000, 168'h000000000000140005000000000000000000000000, 168'h000000000000200000001000000000000000000000, 168'h000000000000404000000000000000000000000000, 168'h000000000000810000000000000000000000000102, 168'h000000000001000040000000000000000000000000, 168'h000000000003000000000000006000000000000000, 168'h000000000005000000000000000000000000000000, 168'h000000000008000000004000000000000000000000, 168'h000000000018000000000000000000000000030000, 168'h000000000030000000030000000000000000000000, 168'h000000000060000000000000000000000000000000, 168'h0000000000a0000014000000000000000000000000, 168'h000000000108000000000000000000000000000000, 168'h000000000240000000000000000000000000000000, 168'h000000000600000000000c00000000000000000000, 168'h000000000800000040000000000000000000000000, 168'h000000001800000000000300000000000000000000, 168'h000000002000000000000010000000000000000000, 168'h000000004008000000000000000000000000000000, 168'h00000000c000000000000000000000000000000600, 168'h000000010000080000000000000000000000000000, 168'h000000030600000000000000000000000000000000, 168'h00000004a400000000000000000000000000000000, 168'h000000080000004000000000000000000000000000, 168'h000000180000003000000000000000000000000000, 168'h000000200001000000000000000000000000000000, 168'h000000600006000000000000000000000000000000, 168'h000000c00000000000000006000000000000000000, 168'h000001000000000000100000000000000000000000, 168'h000003000000000000006000000000000000000000, 168'h000006000000003000000000000000000000000000, 168'h000008000001000000000000000000000000000000, 168'h00001800000000000000000000000000c000000000, 168'h000020000000000001000000000000000000000000, 168'h000048000000000000000000000000000000000000, 168'h0000c0000000000000006000000000000000000000, 168'h000180000000000000000000000000000000000000, 168'h000280000000000000000000000000000005000000, 168'h00060000000c000000000000000000000000000000, 168'h000c00000000000000000000000000018000000000, 168'h001800000600000000000000000000000000000000, 168'h003000000c00000000000000000000000000000000, 168'h004000000080000000000000000000000000000000, 168'h00c000300000000000000000000000000000000000, 168'h010000400000000000000000000000000000000000, 168'h030000000000000000000006000000000000000000, 168'h0600000000000000c0000000000000000000000000, 168'h0c0060000000000000000000000000000000000000, 168'h180000006000000000000000000000000000000000, 168'h3000000000c0000000000000000000000000000000, 168'h410000000000000000000000000000000000000000, 168'ha00140000000000000000000000000000000000000};
	wire lockup;
	wire [LfsrDw - 1:0] lfsr_d;
	reg [LfsrDw - 1:0] lfsr_q;
	wire [LfsrDw - 1:0] next_lfsr_state;
	wire [LfsrDw - 1:0] coeffs;
	generate
		function automatic [63:0] sv2v_cast_64;
			input reg [63:0] inp;
			sv2v_cast_64 = inp;
		endfunction
		if (sv2v_cast_64(LfsrType) == sv2v_cast_64("GAL_XOR")) begin : gen_gal_xor
			if (CustomCoeffs > 0) begin : gen_custom
				assign coeffs = CustomCoeffs[LfsrDw - 1:0];
			end
			else begin : gen_lut
				assign coeffs = GAL_XOR_COEFFS[((60 - (LfsrDw - GAL_XOR_LUT_OFF)) * 64) + (LfsrDw - 1)-:LfsrDw];
			end
			function automatic [LfsrDw - 1:0] sv2v_cast_FFBD2;
				input reg [LfsrDw - 1:0] inp;
				sv2v_cast_FFBD2 = inp;
			endfunction
			assign next_lfsr_state = (sv2v_cast_FFBD2(entropy_i) ^ ({LfsrDw {lfsr_q[0]}} & coeffs)) ^ (lfsr_q >> 1);
			assign lockup = ~(|lfsr_q);
		end
		else begin
			function automatic [63:0] sv2v_cast_64;
				input reg [63:0] inp;
				sv2v_cast_64 = inp;
			endfunction
			if (sv2v_cast_64(LfsrType) == "FIB_XNOR") begin : gen_fib_xnor
				if (CustomCoeffs > 0) begin : gen_custom
					assign coeffs = CustomCoeffs[LfsrDw - 1:0];
				end
				else begin : gen_lut
					assign coeffs = FIB_XNOR_COEFFS[((165 - (LfsrDw - FIB_XNOR_LUT_OFF)) * 168) + (LfsrDw - 1)-:LfsrDw];
				end
				function automatic [LfsrDw - 1:0] sv2v_cast_FFBD2;
					input reg [LfsrDw - 1:0] inp;
					sv2v_cast_FFBD2 = inp;
				endfunction
				assign next_lfsr_state = sv2v_cast_FFBD2(entropy_i) ^ {lfsr_q[LfsrDw - 2:0], ~(^(lfsr_q & coeffs))};
				assign lockup = &lfsr_q;
			end
		end
	endgenerate
	assign lfsr_d = (seed_en_i ? seed_i : (lfsr_en_i && lockup ? DefaultSeed : (lfsr_en_i ? next_lfsr_state : lfsr_q)));
	assign state_o = lfsr_q[StateOutDw - 1:0];
	always @(posedge clk_i or negedge rst_ni) begin : p_reg
		if (!rst_ni)
			lfsr_q <= DefaultSeed;
		else
			lfsr_q <= lfsr_d;
	end
endmodule
