VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spm
  CLASS BLOCK ;
  FOREIGN spm ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.680 BY 131.400 ;
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.850 127.400 95.130 131.400 ;
    END
  END clk
  PIN p
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END p
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END rst
  PIN x[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END x[0]
  PIN x[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END x[10]
  PIN x[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END x[11]
  PIN x[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 116.680 13.640 120.680 14.240 ;
    END
  END x[12]
  PIN x[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END x[13]
  PIN x[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 127.400 50.970 131.400 ;
    END
  END x[14]
  PIN x[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 127.400 17.850 131.400 ;
    END
  END x[15]
  PIN x[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 127.400 73.050 131.400 ;
    END
  END x[16]
  PIN x[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END x[17]
  PIN x[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 116.680 29.960 120.680 30.560 ;
    END
  END x[18]
  PIN x[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END x[19]
  PIN x[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END x[1]
  PIN x[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END x[20]
  PIN x[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 116.680 111.560 120.680 112.160 ;
    END
  END x[21]
  PIN x[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END x[22]
  PIN x[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.890 127.400 106.170 131.400 ;
    END
  END x[23]
  PIN x[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.650 127.400 39.930 131.400 ;
    END
  END x[24]
  PIN x[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 116.680 95.240 120.680 95.840 ;
    END
  END x[25]
  PIN x[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END x[26]
  PIN x[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END x[27]
  PIN x[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 116.680 78.920 120.680 79.520 ;
    END
  END x[28]
  PIN x[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END x[29]
  PIN x[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END x[2]
  PIN x[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 116.680 46.280 120.680 46.880 ;
    END
  END x[30]
  PIN x[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 116.680 62.600 120.680 63.200 ;
    END
  END x[31]
  PIN x[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.530 127.400 6.810 131.400 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.810 127.400 84.090 131.400 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 127.400 62.010 131.400 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END x[7]
  PIN x[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 127.400 28.890 131.400 ;
    END
  END x[8]
  PIN x[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.930 127.400 117.210 131.400 ;
    END
  END x[9]
  PIN y
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END y
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.965 10.640 24.565 119.920 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 41.215 10.640 42.815 119.920 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 115.000 119.765 ;
      LAYER met1 ;
        RECT 2.830 10.640 115.000 120.320 ;
      LAYER met2 ;
        RECT 2.860 127.120 6.250 127.400 ;
        RECT 7.090 127.120 17.290 127.400 ;
        RECT 18.130 127.120 28.330 127.400 ;
        RECT 29.170 127.120 39.370 127.400 ;
        RECT 40.210 127.120 50.410 127.400 ;
        RECT 51.250 127.120 61.450 127.400 ;
        RECT 62.290 127.120 72.490 127.400 ;
        RECT 73.330 127.120 83.530 127.400 ;
        RECT 84.370 127.120 94.570 127.400 ;
        RECT 95.410 127.120 105.610 127.400 ;
        RECT 106.450 127.120 116.650 127.400 ;
        RECT 2.860 4.280 117.210 127.120 ;
        RECT 3.410 4.000 13.610 4.280 ;
        RECT 14.450 4.000 24.650 4.280 ;
        RECT 25.490 4.000 35.690 4.280 ;
        RECT 36.530 4.000 46.730 4.280 ;
        RECT 47.570 4.000 57.770 4.280 ;
        RECT 58.610 4.000 68.810 4.280 ;
        RECT 69.650 4.000 79.850 4.280 ;
        RECT 80.690 4.000 90.890 4.280 ;
        RECT 91.730 4.000 101.930 4.280 ;
        RECT 102.770 4.000 112.970 4.280 ;
        RECT 113.810 4.000 117.210 4.280 ;
      LAYER met3 ;
        RECT 4.000 118.000 117.235 119.845 ;
        RECT 4.400 116.600 117.235 118.000 ;
        RECT 4.000 112.560 117.235 116.600 ;
        RECT 4.000 111.160 116.280 112.560 ;
        RECT 4.000 101.680 117.235 111.160 ;
        RECT 4.400 100.280 117.235 101.680 ;
        RECT 4.000 96.240 117.235 100.280 ;
        RECT 4.000 94.840 116.280 96.240 ;
        RECT 4.000 85.360 117.235 94.840 ;
        RECT 4.400 83.960 117.235 85.360 ;
        RECT 4.000 79.920 117.235 83.960 ;
        RECT 4.000 78.520 116.280 79.920 ;
        RECT 4.000 69.040 117.235 78.520 ;
        RECT 4.400 67.640 117.235 69.040 ;
        RECT 4.000 63.600 117.235 67.640 ;
        RECT 4.000 62.200 116.280 63.600 ;
        RECT 4.000 52.720 117.235 62.200 ;
        RECT 4.400 51.320 117.235 52.720 ;
        RECT 4.000 47.280 117.235 51.320 ;
        RECT 4.000 45.880 116.280 47.280 ;
        RECT 4.000 36.400 117.235 45.880 ;
        RECT 4.400 35.000 117.235 36.400 ;
        RECT 4.000 30.960 117.235 35.000 ;
        RECT 4.000 29.560 116.280 30.960 ;
        RECT 4.000 20.080 117.235 29.560 ;
        RECT 4.400 18.680 117.235 20.080 ;
        RECT 4.000 14.640 117.235 18.680 ;
        RECT 4.000 13.240 116.280 14.640 ;
        RECT 4.000 10.715 117.235 13.240 ;
      LAYER met4 ;
        RECT 43.215 10.640 97.550 119.920 ;
  END
END spm
END LIBRARY

