//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[22][0]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Tue Feb 25 16:43:51 2020
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

`include "../fpga_defines.v"
// ----- Verilog module for sb_22__0_ -----
module sb_22__0_(pReset,
                 prog_clk,
                 chany_top_in_1_,
                 chany_top_in_3_,
                 chany_top_in_5_,
                 chany_top_in_7_,
                 chany_top_in_9_,
                 chany_top_in_11_,
                 chany_top_in_13_,
                 chany_top_in_15_,
                 chany_top_in_17_,
                 chany_top_in_19_,
                 chany_top_in_21_,
                 chany_top_in_23_,
                 chany_top_in_25_,
                 chany_top_in_27_,
                 chany_top_in_29_,
                 chany_top_in_31_,
                 chany_top_in_33_,
                 chany_top_in_35_,
                 chany_top_in_37_,
                 chany_top_in_39_,
                 chany_top_in_41_,
                 chany_top_in_43_,
                 chany_top_in_45_,
                 chany_top_in_47_,
                 chany_top_in_49_,
                 chany_top_in_51_,
                 chany_top_in_53_,
                 chany_top_in_55_,
                 chany_top_in_57_,
                 chany_top_in_59_,
                 chany_top_in_61_,
                 chany_top_in_63_,
                 chany_top_in_65_,
                 chany_top_in_67_,
                 chany_top_in_69_,
                 chany_top_in_71_,
                 chany_top_in_73_,
                 chany_top_in_75_,
                 chany_top_in_77_,
                 chany_top_in_79_,
                 chany_top_in_81_,
                 chany_top_in_83_,
                 chany_top_in_85_,
                 chany_top_in_87_,
                 chany_top_in_89_,
                 chany_top_in_91_,
                 chany_top_in_93_,
                 chany_top_in_95_,
                 chany_top_in_97_,
                 chany_top_in_99_,
                 chany_top_in_101_,
                 chany_top_in_103_,
                 chany_top_in_105_,
                 chany_top_in_107_,
                 chany_top_in_109_,
                 chany_top_in_111_,
                 chany_top_in_113_,
                 chany_top_in_115_,
                 chany_top_in_117_,
                 chany_top_in_119_,
                 top_left_grid_pin_30_,
                 top_left_grid_pin_31_,
                 top_left_grid_pin_32_,
                 top_left_grid_pin_33_,
                 top_left_grid_pin_34_,
                 top_right_grid_pin_1_,
                 chanx_left_in_0_,
                 chanx_left_in_2_,
                 chanx_left_in_4_,
                 chanx_left_in_6_,
                 chanx_left_in_8_,
                 chanx_left_in_10_,
                 chanx_left_in_12_,
                 chanx_left_in_14_,
                 chanx_left_in_16_,
                 chanx_left_in_18_,
                 chanx_left_in_20_,
                 chanx_left_in_22_,
                 chanx_left_in_24_,
                 chanx_left_in_26_,
                 chanx_left_in_28_,
                 chanx_left_in_30_,
                 chanx_left_in_32_,
                 chanx_left_in_34_,
                 chanx_left_in_36_,
                 chanx_left_in_38_,
                 chanx_left_in_40_,
                 chanx_left_in_42_,
                 chanx_left_in_44_,
                 chanx_left_in_46_,
                 chanx_left_in_48_,
                 chanx_left_in_50_,
                 chanx_left_in_52_,
                 chanx_left_in_54_,
                 chanx_left_in_56_,
                 chanx_left_in_58_,
                 chanx_left_in_60_,
                 chanx_left_in_62_,
                 chanx_left_in_64_,
                 chanx_left_in_66_,
                 chanx_left_in_68_,
                 chanx_left_in_70_,
                 chanx_left_in_72_,
                 chanx_left_in_74_,
                 chanx_left_in_76_,
                 chanx_left_in_78_,
                 chanx_left_in_80_,
                 chanx_left_in_82_,
                 chanx_left_in_84_,
                 chanx_left_in_86_,
                 chanx_left_in_88_,
                 chanx_left_in_90_,
                 chanx_left_in_92_,
                 chanx_left_in_94_,
                 chanx_left_in_96_,
                 chanx_left_in_98_,
                 chanx_left_in_100_,
                 chanx_left_in_102_,
                 chanx_left_in_104_,
                 chanx_left_in_106_,
                 chanx_left_in_108_,
                 chanx_left_in_110_,
                 chanx_left_in_112_,
                 chanx_left_in_114_,
                 chanx_left_in_116_,
                 chanx_left_in_118_,
                 left_top_grid_pin_35_,
                 left_top_grid_pin_36_,
                 left_top_grid_pin_37_,
                 left_top_grid_pin_38_,
                 left_top_grid_pin_39_,
                 left_bottom_grid_pin_1_,
                 ccff_head,
                 chany_top_out_0_,
                 chany_top_out_2_,
                 chany_top_out_4_,
                 chany_top_out_6_,
                 chany_top_out_8_,
                 chany_top_out_10_,
                 chany_top_out_12_,
                 chany_top_out_14_,
                 chany_top_out_16_,
                 chany_top_out_18_,
                 chany_top_out_20_,
                 chany_top_out_22_,
                 chany_top_out_24_,
                 chany_top_out_26_,
                 chany_top_out_28_,
                 chany_top_out_30_,
                 chany_top_out_32_,
                 chany_top_out_34_,
                 chany_top_out_36_,
                 chany_top_out_38_,
                 chany_top_out_40_,
                 chany_top_out_42_,
                 chany_top_out_44_,
                 chany_top_out_46_,
                 chany_top_out_48_,
                 chany_top_out_50_,
                 chany_top_out_52_,
                 chany_top_out_54_,
                 chany_top_out_56_,
                 chany_top_out_58_,
                 chany_top_out_60_,
                 chany_top_out_62_,
                 chany_top_out_64_,
                 chany_top_out_66_,
                 chany_top_out_68_,
                 chany_top_out_70_,
                 chany_top_out_72_,
                 chany_top_out_74_,
                 chany_top_out_76_,
                 chany_top_out_78_,
                 chany_top_out_80_,
                 chany_top_out_82_,
                 chany_top_out_84_,
                 chany_top_out_86_,
                 chany_top_out_88_,
                 chany_top_out_90_,
                 chany_top_out_92_,
                 chany_top_out_94_,
                 chany_top_out_96_,
                 chany_top_out_98_,
                 chany_top_out_100_,
                 chany_top_out_102_,
                 chany_top_out_104_,
                 chany_top_out_106_,
                 chany_top_out_108_,
                 chany_top_out_110_,
                 chany_top_out_112_,
                 chany_top_out_114_,
                 chany_top_out_116_,
                 chany_top_out_118_,
                 chanx_left_out_1_,
                 chanx_left_out_3_,
                 chanx_left_out_5_,
                 chanx_left_out_7_,
                 chanx_left_out_9_,
                 chanx_left_out_11_,
                 chanx_left_out_13_,
                 chanx_left_out_15_,
                 chanx_left_out_17_,
                 chanx_left_out_19_,
                 chanx_left_out_21_,
                 chanx_left_out_23_,
                 chanx_left_out_25_,
                 chanx_left_out_27_,
                 chanx_left_out_29_,
                 chanx_left_out_31_,
                 chanx_left_out_33_,
                 chanx_left_out_35_,
                 chanx_left_out_37_,
                 chanx_left_out_39_,
                 chanx_left_out_41_,
                 chanx_left_out_43_,
                 chanx_left_out_45_,
                 chanx_left_out_47_,
                 chanx_left_out_49_,
                 chanx_left_out_51_,
                 chanx_left_out_53_,
                 chanx_left_out_55_,
                 chanx_left_out_57_,
                 chanx_left_out_59_,
                 chanx_left_out_61_,
                 chanx_left_out_63_,
                 chanx_left_out_65_,
                 chanx_left_out_67_,
                 chanx_left_out_69_,
                 chanx_left_out_71_,
                 chanx_left_out_73_,
                 chanx_left_out_75_,
                 chanx_left_out_77_,
                 chanx_left_out_79_,
                 chanx_left_out_81_,
                 chanx_left_out_83_,
                 chanx_left_out_85_,
                 chanx_left_out_87_,
                 chanx_left_out_89_,
                 chanx_left_out_91_,
                 chanx_left_out_93_,
                 chanx_left_out_95_,
                 chanx_left_out_97_,
                 chanx_left_out_99_,
                 chanx_left_out_101_,
                 chanx_left_out_103_,
                 chanx_left_out_105_,
                 chanx_left_out_107_,
                 chanx_left_out_109_,
                 chanx_left_out_111_,
                 chanx_left_out_113_,
                 chanx_left_out_115_,
                 chanx_left_out_117_,
                 chanx_left_out_119_,
                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] chany_top_in_1_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_3_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_5_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_7_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_9_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_11_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_13_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_15_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_17_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_19_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_21_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_23_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_25_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_27_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_29_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_31_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_33_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_35_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_37_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_39_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_41_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_43_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_45_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_47_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_49_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_51_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_53_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_55_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_57_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_59_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_61_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_63_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_65_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_67_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_69_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_71_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_73_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_75_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_77_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_79_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_81_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_83_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_85_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_87_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_89_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_91_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_93_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_95_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_97_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_99_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_101_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_103_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_105_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_107_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_109_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_111_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_113_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_115_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_117_;
//----- INPUT PORTS -----
input [0:0] chany_top_in_119_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_pin_30_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_pin_31_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_pin_32_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_pin_33_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_pin_34_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_pin_1_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_0_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_2_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_4_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_6_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_8_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_10_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_12_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_14_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_16_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_18_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_20_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_22_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_24_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_26_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_28_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_30_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_32_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_34_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_36_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_38_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_40_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_42_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_44_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_46_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_48_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_50_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_52_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_54_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_56_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_58_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_60_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_62_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_64_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_66_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_68_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_70_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_72_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_74_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_76_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_78_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_80_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_82_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_84_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_86_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_88_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_90_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_92_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_94_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_96_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_98_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_100_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_102_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_104_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_106_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_108_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_110_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_112_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_114_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_116_;
//----- INPUT PORTS -----
input [0:0] chanx_left_in_118_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_pin_35_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_pin_36_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_pin_37_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_pin_38_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_pin_39_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_pin_1_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_0_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_2_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_4_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_6_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_8_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_10_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_12_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_14_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_16_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_18_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_20_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_22_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_24_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_26_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_28_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_30_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_32_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_34_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_36_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_38_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_40_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_42_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_44_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_46_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_48_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_50_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_52_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_54_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_56_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_58_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_60_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_62_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_64_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_66_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_68_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_70_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_72_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_74_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_76_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_78_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_80_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_82_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_84_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_86_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_88_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_90_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_92_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_94_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_96_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_98_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_100_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_102_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_104_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_106_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_108_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_110_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_112_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_114_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_116_;
//----- OUTPUT PORTS -----
output [0:0] chany_top_out_118_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_1_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_3_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_5_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_7_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_9_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_11_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_13_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_15_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_17_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_19_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_21_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_23_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_25_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_27_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_29_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_31_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_33_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_35_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_37_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_39_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_41_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_43_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_45_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_47_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_49_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_51_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_53_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_55_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_57_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_59_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_61_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_63_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_65_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_67_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_69_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_71_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_73_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_75_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_77_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_79_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_81_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_83_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_85_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_87_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_89_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_91_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_93_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_95_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_97_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_99_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_101_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_103_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_105_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_107_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_109_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_111_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_113_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_115_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_117_;
//----- OUTPUT PORTS -----
output [0:0] chanx_left_out_119_;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_like_tapbuf_size2_0_sram;
wire [0:1] mux_tree_like_tapbuf_size2_0_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_10_sram;
wire [0:1] mux_tree_like_tapbuf_size2_10_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_11_sram;
wire [0:1] mux_tree_like_tapbuf_size2_11_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_12_sram;
wire [0:1] mux_tree_like_tapbuf_size2_12_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_13_sram;
wire [0:1] mux_tree_like_tapbuf_size2_13_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_14_sram;
wire [0:1] mux_tree_like_tapbuf_size2_14_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_15_sram;
wire [0:1] mux_tree_like_tapbuf_size2_15_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_16_sram;
wire [0:1] mux_tree_like_tapbuf_size2_16_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_17_sram;
wire [0:1] mux_tree_like_tapbuf_size2_17_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_18_sram;
wire [0:1] mux_tree_like_tapbuf_size2_18_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_19_sram;
wire [0:1] mux_tree_like_tapbuf_size2_19_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_1_sram;
wire [0:1] mux_tree_like_tapbuf_size2_1_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_20_sram;
wire [0:1] mux_tree_like_tapbuf_size2_20_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_21_sram;
wire [0:1] mux_tree_like_tapbuf_size2_21_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_22_sram;
wire [0:1] mux_tree_like_tapbuf_size2_22_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_23_sram;
wire [0:1] mux_tree_like_tapbuf_size2_23_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_24_sram;
wire [0:1] mux_tree_like_tapbuf_size2_24_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_25_sram;
wire [0:1] mux_tree_like_tapbuf_size2_25_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_26_sram;
wire [0:1] mux_tree_like_tapbuf_size2_26_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_27_sram;
wire [0:1] mux_tree_like_tapbuf_size2_27_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_28_sram;
wire [0:1] mux_tree_like_tapbuf_size2_28_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_29_sram;
wire [0:1] mux_tree_like_tapbuf_size2_29_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_2_sram;
wire [0:1] mux_tree_like_tapbuf_size2_2_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_30_sram;
wire [0:1] mux_tree_like_tapbuf_size2_30_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_31_sram;
wire [0:1] mux_tree_like_tapbuf_size2_31_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_32_sram;
wire [0:1] mux_tree_like_tapbuf_size2_32_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_33_sram;
wire [0:1] mux_tree_like_tapbuf_size2_33_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_34_sram;
wire [0:1] mux_tree_like_tapbuf_size2_34_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_35_sram;
wire [0:1] mux_tree_like_tapbuf_size2_35_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_36_sram;
wire [0:1] mux_tree_like_tapbuf_size2_36_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_37_sram;
wire [0:1] mux_tree_like_tapbuf_size2_37_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_38_sram;
wire [0:1] mux_tree_like_tapbuf_size2_38_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_39_sram;
wire [0:1] mux_tree_like_tapbuf_size2_39_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_3_sram;
wire [0:1] mux_tree_like_tapbuf_size2_3_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_40_sram;
wire [0:1] mux_tree_like_tapbuf_size2_40_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_41_sram;
wire [0:1] mux_tree_like_tapbuf_size2_41_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_42_sram;
wire [0:1] mux_tree_like_tapbuf_size2_42_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_43_sram;
wire [0:1] mux_tree_like_tapbuf_size2_43_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_44_sram;
wire [0:1] mux_tree_like_tapbuf_size2_44_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_45_sram;
wire [0:1] mux_tree_like_tapbuf_size2_45_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_46_sram;
wire [0:1] mux_tree_like_tapbuf_size2_46_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_47_sram;
wire [0:1] mux_tree_like_tapbuf_size2_47_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_48_sram;
wire [0:1] mux_tree_like_tapbuf_size2_48_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_49_sram;
wire [0:1] mux_tree_like_tapbuf_size2_49_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_4_sram;
wire [0:1] mux_tree_like_tapbuf_size2_4_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_50_sram;
wire [0:1] mux_tree_like_tapbuf_size2_50_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_51_sram;
wire [0:1] mux_tree_like_tapbuf_size2_51_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_52_sram;
wire [0:1] mux_tree_like_tapbuf_size2_52_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_53_sram;
wire [0:1] mux_tree_like_tapbuf_size2_53_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_54_sram;
wire [0:1] mux_tree_like_tapbuf_size2_54_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_55_sram;
wire [0:1] mux_tree_like_tapbuf_size2_55_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_56_sram;
wire [0:1] mux_tree_like_tapbuf_size2_56_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_57_sram;
wire [0:1] mux_tree_like_tapbuf_size2_57_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_58_sram;
wire [0:1] mux_tree_like_tapbuf_size2_58_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_59_sram;
wire [0:1] mux_tree_like_tapbuf_size2_59_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_5_sram;
wire [0:1] mux_tree_like_tapbuf_size2_5_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_60_sram;
wire [0:1] mux_tree_like_tapbuf_size2_60_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_61_sram;
wire [0:1] mux_tree_like_tapbuf_size2_61_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_62_sram;
wire [0:1] mux_tree_like_tapbuf_size2_62_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_63_sram;
wire [0:1] mux_tree_like_tapbuf_size2_63_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_64_sram;
wire [0:1] mux_tree_like_tapbuf_size2_64_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_65_sram;
wire [0:1] mux_tree_like_tapbuf_size2_65_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_66_sram;
wire [0:1] mux_tree_like_tapbuf_size2_66_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_67_sram;
wire [0:1] mux_tree_like_tapbuf_size2_67_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_68_sram;
wire [0:1] mux_tree_like_tapbuf_size2_68_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_69_sram;
wire [0:1] mux_tree_like_tapbuf_size2_69_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_6_sram;
wire [0:1] mux_tree_like_tapbuf_size2_6_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_70_sram;
wire [0:1] mux_tree_like_tapbuf_size2_70_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_71_sram;
wire [0:1] mux_tree_like_tapbuf_size2_71_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_72_sram;
wire [0:1] mux_tree_like_tapbuf_size2_72_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_73_sram;
wire [0:1] mux_tree_like_tapbuf_size2_73_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_74_sram;
wire [0:1] mux_tree_like_tapbuf_size2_74_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_75_sram;
wire [0:1] mux_tree_like_tapbuf_size2_75_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_76_sram;
wire [0:1] mux_tree_like_tapbuf_size2_76_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_77_sram;
wire [0:1] mux_tree_like_tapbuf_size2_77_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_78_sram;
wire [0:1] mux_tree_like_tapbuf_size2_78_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_79_sram;
wire [0:1] mux_tree_like_tapbuf_size2_79_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_7_sram;
wire [0:1] mux_tree_like_tapbuf_size2_7_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_80_sram;
wire [0:1] mux_tree_like_tapbuf_size2_80_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_81_sram;
wire [0:1] mux_tree_like_tapbuf_size2_81_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_82_sram;
wire [0:1] mux_tree_like_tapbuf_size2_82_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_83_sram;
wire [0:1] mux_tree_like_tapbuf_size2_83_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_84_sram;
wire [0:1] mux_tree_like_tapbuf_size2_84_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_85_sram;
wire [0:1] mux_tree_like_tapbuf_size2_85_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_86_sram;
wire [0:1] mux_tree_like_tapbuf_size2_86_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_87_sram;
wire [0:1] mux_tree_like_tapbuf_size2_87_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_8_sram;
wire [0:1] mux_tree_like_tapbuf_size2_8_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size2_9_sram;
wire [0:1] mux_tree_like_tapbuf_size2_9_sram_inv;
wire [0:0] mux_tree_like_tapbuf_size2_mem_0_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_10_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_11_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_12_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_13_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_14_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_15_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_16_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_17_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_18_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_19_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_1_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_20_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_21_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_22_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_23_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_24_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_25_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_26_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_27_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_28_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_29_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_2_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_30_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_31_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_32_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_33_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_34_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_35_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_36_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_37_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_38_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_39_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_3_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_40_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_41_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_42_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_43_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_44_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_45_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_46_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_47_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_48_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_49_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_4_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_50_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_51_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_52_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_53_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_54_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_55_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_56_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_57_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_58_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_59_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_5_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_60_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_61_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_62_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_63_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_64_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_65_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_66_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_67_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_68_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_69_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_6_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_70_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_71_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_72_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_73_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_74_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_75_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_76_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_77_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_78_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_79_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_7_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_80_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_81_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_82_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_83_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_84_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_85_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_86_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_8_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size2_mem_9_ccff_tail;
wire [0:1] mux_tree_like_tapbuf_size3_0_sram;
wire [0:1] mux_tree_like_tapbuf_size3_0_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size3_1_sram;
wire [0:1] mux_tree_like_tapbuf_size3_1_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size3_2_sram;
wire [0:1] mux_tree_like_tapbuf_size3_2_sram_inv;
wire [0:1] mux_tree_like_tapbuf_size3_3_sram;
wire [0:1] mux_tree_like_tapbuf_size3_3_sram_inv;
wire [0:0] mux_tree_like_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_tree_like_tapbuf_size3_mem_3_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out_111_[0] = chany_top_in_11_[0];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out_109_[0] = chany_top_in_13_[0];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out_95_[0] = chany_top_in_27_[0];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out_93_[0] = chany_top_in_29_[0];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out_79_[0] = chany_top_in_43_[0];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out_77_[0] = chany_top_in_45_[0];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out_63_[0] = chany_top_in_59_[0];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out_61_[0] = chany_top_in_61_[0];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out_47_[0] = chany_top_in_75_[0];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out_45_[0] = chany_top_in_77_[0];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out_31_[0] = chany_top_in_91_[0];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out_29_[0] = chany_top_in_93_[0];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out_15_[0] = chany_top_in_107_[0];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_left_out_13_[0] = chany_top_in_109_[0];
// ----- Local connection due to Wire 71 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out_110_[0] = chanx_left_in_10_[0];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out_108_[0] = chanx_left_in_12_[0];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out_94_[0] = chanx_left_in_26_[0];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out_92_[0] = chanx_left_in_28_[0];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out_78_[0] = chanx_left_in_42_[0];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out_76_[0] = chanx_left_in_44_[0];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out_62_[0] = chanx_left_in_58_[0];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out_60_[0] = chanx_left_in_60_[0];
// ----- Local connection due to Wire 103 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out_46_[0] = chanx_left_in_74_[0];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out_44_[0] = chanx_left_in_76_[0];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out_30_[0] = chanx_left_in_90_[0];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out_28_[0] = chanx_left_in_92_[0];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out_14_[0] = chanx_left_in_106_[0];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out_12_[0] = chanx_left_in_108_[0];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_like_tapbuf_size2 mux_top_track_0 (
		.in({top_left_grid_pin_30_[0], chanx_left_in_0_[0]}),
		.sram(mux_tree_like_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_0_sram_inv[0:1]),
		.out(chany_top_out_0_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_2 (
		.in({top_left_grid_pin_31_[0], chanx_left_in_118_[0]}),
		.sram(mux_tree_like_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_1_sram_inv[0:1]),
		.out(chany_top_out_2_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_4 (
		.in({top_left_grid_pin_32_[0], chanx_left_in_116_[0]}),
		.sram(mux_tree_like_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_2_sram_inv[0:1]),
		.out(chany_top_out_4_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_6 (
		.in({top_left_grid_pin_33_[0], chanx_left_in_114_[0]}),
		.sram(mux_tree_like_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_3_sram_inv[0:1]),
		.out(chany_top_out_6_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_8 (
		.in({top_left_grid_pin_34_[0], chanx_left_in_112_[0]}),
		.sram(mux_tree_like_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_4_sram_inv[0:1]),
		.out(chany_top_out_8_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_10 (
		.in({top_right_grid_pin_1_[0], chanx_left_in_110_[0]}),
		.sram(mux_tree_like_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_5_sram_inv[0:1]),
		.out(chany_top_out_10_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_20 (
		.in({top_left_grid_pin_32_[0], chanx_left_in_100_[0]}),
		.sram(mux_tree_like_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_6_sram_inv[0:1]),
		.out(chany_top_out_20_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_22 (
		.in({top_left_grid_pin_33_[0], chanx_left_in_98_[0]}),
		.sram(mux_tree_like_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_7_sram_inv[0:1]),
		.out(chany_top_out_22_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_24 (
		.in({top_left_grid_pin_34_[0], chanx_left_in_96_[0]}),
		.sram(mux_tree_like_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_8_sram_inv[0:1]),
		.out(chany_top_out_24_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_26 (
		.in({top_right_grid_pin_1_[0], chanx_left_in_94_[0]}),
		.sram(mux_tree_like_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_9_sram_inv[0:1]),
		.out(chany_top_out_26_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_32 (
		.in({top_left_grid_pin_30_[0], chanx_left_in_88_[0]}),
		.sram(mux_tree_like_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_10_sram_inv[0:1]),
		.out(chany_top_out_32_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_34 (
		.in({top_left_grid_pin_31_[0], chanx_left_in_86_[0]}),
		.sram(mux_tree_like_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_11_sram_inv[0:1]),
		.out(chany_top_out_34_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_36 (
		.in({top_left_grid_pin_32_[0], chanx_left_in_84_[0]}),
		.sram(mux_tree_like_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_12_sram_inv[0:1]),
		.out(chany_top_out_36_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_38 (
		.in({top_left_grid_pin_33_[0], chanx_left_in_82_[0]}),
		.sram(mux_tree_like_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_13_sram_inv[0:1]),
		.out(chany_top_out_38_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_40 (
		.in({top_left_grid_pin_34_[0], chanx_left_in_80_[0]}),
		.sram(mux_tree_like_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_14_sram_inv[0:1]),
		.out(chany_top_out_40_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_42 (
		.in({top_right_grid_pin_1_[0], chanx_left_in_78_[0]}),
		.sram(mux_tree_like_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_15_sram_inv[0:1]),
		.out(chany_top_out_42_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_48 (
		.in({top_left_grid_pin_30_[0], chanx_left_in_72_[0]}),
		.sram(mux_tree_like_tapbuf_size2_16_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_16_sram_inv[0:1]),
		.out(chany_top_out_48_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_50 (
		.in({top_left_grid_pin_31_[0], chanx_left_in_70_[0]}),
		.sram(mux_tree_like_tapbuf_size2_17_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_17_sram_inv[0:1]),
		.out(chany_top_out_50_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_52 (
		.in({top_left_grid_pin_32_[0], chanx_left_in_68_[0]}),
		.sram(mux_tree_like_tapbuf_size2_18_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_18_sram_inv[0:1]),
		.out(chany_top_out_52_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_54 (
		.in({top_left_grid_pin_33_[0], chanx_left_in_66_[0]}),
		.sram(mux_tree_like_tapbuf_size2_19_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_19_sram_inv[0:1]),
		.out(chany_top_out_54_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_56 (
		.in({top_left_grid_pin_34_[0], chanx_left_in_64_[0]}),
		.sram(mux_tree_like_tapbuf_size2_20_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_20_sram_inv[0:1]),
		.out(chany_top_out_56_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_58 (
		.in({top_right_grid_pin_1_[0], chanx_left_in_62_[0]}),
		.sram(mux_tree_like_tapbuf_size2_21_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_21_sram_inv[0:1]),
		.out(chany_top_out_58_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_64 (
		.in({top_left_grid_pin_30_[0], chanx_left_in_56_[0]}),
		.sram(mux_tree_like_tapbuf_size2_22_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_22_sram_inv[0:1]),
		.out(chany_top_out_64_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_66 (
		.in({top_left_grid_pin_31_[0], chanx_left_in_54_[0]}),
		.sram(mux_tree_like_tapbuf_size2_23_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_23_sram_inv[0:1]),
		.out(chany_top_out_66_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_68 (
		.in({top_left_grid_pin_32_[0], chanx_left_in_52_[0]}),
		.sram(mux_tree_like_tapbuf_size2_24_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_24_sram_inv[0:1]),
		.out(chany_top_out_68_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_70 (
		.in({top_left_grid_pin_33_[0], chanx_left_in_50_[0]}),
		.sram(mux_tree_like_tapbuf_size2_25_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_25_sram_inv[0:1]),
		.out(chany_top_out_70_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_72 (
		.in({top_left_grid_pin_34_[0], chanx_left_in_48_[0]}),
		.sram(mux_tree_like_tapbuf_size2_26_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_26_sram_inv[0:1]),
		.out(chany_top_out_72_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_74 (
		.in({top_right_grid_pin_1_[0], chanx_left_in_46_[0]}),
		.sram(mux_tree_like_tapbuf_size2_27_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_27_sram_inv[0:1]),
		.out(chany_top_out_74_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_80 (
		.in({top_left_grid_pin_30_[0], chanx_left_in_40_[0]}),
		.sram(mux_tree_like_tapbuf_size2_28_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_28_sram_inv[0:1]),
		.out(chany_top_out_80_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_82 (
		.in({top_left_grid_pin_31_[0], chanx_left_in_38_[0]}),
		.sram(mux_tree_like_tapbuf_size2_29_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_29_sram_inv[0:1]),
		.out(chany_top_out_82_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_84 (
		.in({top_left_grid_pin_32_[0], chanx_left_in_36_[0]}),
		.sram(mux_tree_like_tapbuf_size2_30_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_30_sram_inv[0:1]),
		.out(chany_top_out_84_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_86 (
		.in({top_left_grid_pin_33_[0], chanx_left_in_34_[0]}),
		.sram(mux_tree_like_tapbuf_size2_31_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_31_sram_inv[0:1]),
		.out(chany_top_out_86_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_88 (
		.in({top_left_grid_pin_34_[0], chanx_left_in_32_[0]}),
		.sram(mux_tree_like_tapbuf_size2_32_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_32_sram_inv[0:1]),
		.out(chany_top_out_88_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_90 (
		.in({top_right_grid_pin_1_[0], chanx_left_in_30_[0]}),
		.sram(mux_tree_like_tapbuf_size2_33_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_33_sram_inv[0:1]),
		.out(chany_top_out_90_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_96 (
		.in({top_left_grid_pin_30_[0], chanx_left_in_24_[0]}),
		.sram(mux_tree_like_tapbuf_size2_34_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_34_sram_inv[0:1]),
		.out(chany_top_out_96_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_98 (
		.in({top_left_grid_pin_31_[0], chanx_left_in_22_[0]}),
		.sram(mux_tree_like_tapbuf_size2_35_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_35_sram_inv[0:1]),
		.out(chany_top_out_98_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_100 (
		.in({top_left_grid_pin_32_[0], chanx_left_in_20_[0]}),
		.sram(mux_tree_like_tapbuf_size2_36_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_36_sram_inv[0:1]),
		.out(chany_top_out_100_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_102 (
		.in({top_left_grid_pin_33_[0], chanx_left_in_18_[0]}),
		.sram(mux_tree_like_tapbuf_size2_37_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_37_sram_inv[0:1]),
		.out(chany_top_out_102_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_104 (
		.in({top_left_grid_pin_34_[0], chanx_left_in_16_[0]}),
		.sram(mux_tree_like_tapbuf_size2_38_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_38_sram_inv[0:1]),
		.out(chany_top_out_104_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_106 (
		.in({top_right_grid_pin_1_[0], chanx_left_in_14_[0]}),
		.sram(mux_tree_like_tapbuf_size2_39_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_39_sram_inv[0:1]),
		.out(chany_top_out_106_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_112 (
		.in({top_left_grid_pin_30_[0], chanx_left_in_8_[0]}),
		.sram(mux_tree_like_tapbuf_size2_40_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_40_sram_inv[0:1]),
		.out(chany_top_out_112_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_114 (
		.in({top_left_grid_pin_31_[0], chanx_left_in_6_[0]}),
		.sram(mux_tree_like_tapbuf_size2_41_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_41_sram_inv[0:1]),
		.out(chany_top_out_114_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_116 (
		.in({top_left_grid_pin_32_[0], chanx_left_in_4_[0]}),
		.sram(mux_tree_like_tapbuf_size2_42_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_42_sram_inv[0:1]),
		.out(chany_top_out_116_[0]));

	mux_tree_like_tapbuf_size2 mux_top_track_118 (
		.in({top_left_grid_pin_33_[0], chanx_left_in_2_[0]}),
		.sram(mux_tree_like_tapbuf_size2_43_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_43_sram_inv[0:1]),
		.out(chany_top_out_118_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_1 (
		.in({left_top_grid_pin_35_[0], chany_top_in_1_[0]}),
		.sram(mux_tree_like_tapbuf_size2_44_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_44_sram_inv[0:1]),
		.out(chanx_left_out_1_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_3 (
		.in({left_top_grid_pin_36_[0], chany_top_in_119_[0]}),
		.sram(mux_tree_like_tapbuf_size2_45_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_45_sram_inv[0:1]),
		.out(chanx_left_out_3_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_5 (
		.in({left_top_grid_pin_37_[0], chany_top_in_117_[0]}),
		.sram(mux_tree_like_tapbuf_size2_46_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_46_sram_inv[0:1]),
		.out(chanx_left_out_5_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_7 (
		.in({left_top_grid_pin_38_[0], chany_top_in_115_[0]}),
		.sram(mux_tree_like_tapbuf_size2_47_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_47_sram_inv[0:1]),
		.out(chanx_left_out_7_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_9 (
		.in({left_top_grid_pin_39_[0], chany_top_in_113_[0]}),
		.sram(mux_tree_like_tapbuf_size2_48_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_48_sram_inv[0:1]),
		.out(chanx_left_out_9_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_11 (
		.in({left_bottom_grid_pin_1_[0], chany_top_in_111_[0]}),
		.sram(mux_tree_like_tapbuf_size2_49_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_49_sram_inv[0:1]),
		.out(chanx_left_out_11_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_21 (
		.in({left_top_grid_pin_37_[0], chany_top_in_101_[0]}),
		.sram(mux_tree_like_tapbuf_size2_50_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_50_sram_inv[0:1]),
		.out(chanx_left_out_21_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_23 (
		.in({left_top_grid_pin_38_[0], chany_top_in_99_[0]}),
		.sram(mux_tree_like_tapbuf_size2_51_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_51_sram_inv[0:1]),
		.out(chanx_left_out_23_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_25 (
		.in({left_top_grid_pin_39_[0], chany_top_in_97_[0]}),
		.sram(mux_tree_like_tapbuf_size2_52_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_52_sram_inv[0:1]),
		.out(chanx_left_out_25_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_27 (
		.in({left_bottom_grid_pin_1_[0], chany_top_in_95_[0]}),
		.sram(mux_tree_like_tapbuf_size2_53_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_53_sram_inv[0:1]),
		.out(chanx_left_out_27_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_33 (
		.in({left_top_grid_pin_35_[0], chany_top_in_89_[0]}),
		.sram(mux_tree_like_tapbuf_size2_54_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_54_sram_inv[0:1]),
		.out(chanx_left_out_33_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_35 (
		.in({left_top_grid_pin_36_[0], chany_top_in_87_[0]}),
		.sram(mux_tree_like_tapbuf_size2_55_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_55_sram_inv[0:1]),
		.out(chanx_left_out_35_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_37 (
		.in({left_top_grid_pin_37_[0], chany_top_in_85_[0]}),
		.sram(mux_tree_like_tapbuf_size2_56_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_56_sram_inv[0:1]),
		.out(chanx_left_out_37_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_39 (
		.in({left_top_grid_pin_38_[0], chany_top_in_83_[0]}),
		.sram(mux_tree_like_tapbuf_size2_57_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_57_sram_inv[0:1]),
		.out(chanx_left_out_39_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_41 (
		.in({left_top_grid_pin_39_[0], chany_top_in_81_[0]}),
		.sram(mux_tree_like_tapbuf_size2_58_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_58_sram_inv[0:1]),
		.out(chanx_left_out_41_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_43 (
		.in({left_bottom_grid_pin_1_[0], chany_top_in_79_[0]}),
		.sram(mux_tree_like_tapbuf_size2_59_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_59_sram_inv[0:1]),
		.out(chanx_left_out_43_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_49 (
		.in({left_top_grid_pin_35_[0], chany_top_in_73_[0]}),
		.sram(mux_tree_like_tapbuf_size2_60_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_60_sram_inv[0:1]),
		.out(chanx_left_out_49_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_51 (
		.in({left_top_grid_pin_36_[0], chany_top_in_71_[0]}),
		.sram(mux_tree_like_tapbuf_size2_61_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_61_sram_inv[0:1]),
		.out(chanx_left_out_51_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_53 (
		.in({left_top_grid_pin_37_[0], chany_top_in_69_[0]}),
		.sram(mux_tree_like_tapbuf_size2_62_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_62_sram_inv[0:1]),
		.out(chanx_left_out_53_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_55 (
		.in({left_top_grid_pin_38_[0], chany_top_in_67_[0]}),
		.sram(mux_tree_like_tapbuf_size2_63_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_63_sram_inv[0:1]),
		.out(chanx_left_out_55_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_57 (
		.in({left_top_grid_pin_39_[0], chany_top_in_65_[0]}),
		.sram(mux_tree_like_tapbuf_size2_64_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_64_sram_inv[0:1]),
		.out(chanx_left_out_57_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_59 (
		.in({left_bottom_grid_pin_1_[0], chany_top_in_63_[0]}),
		.sram(mux_tree_like_tapbuf_size2_65_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_65_sram_inv[0:1]),
		.out(chanx_left_out_59_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_65 (
		.in({left_top_grid_pin_35_[0], chany_top_in_57_[0]}),
		.sram(mux_tree_like_tapbuf_size2_66_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_66_sram_inv[0:1]),
		.out(chanx_left_out_65_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_67 (
		.in({left_top_grid_pin_36_[0], chany_top_in_55_[0]}),
		.sram(mux_tree_like_tapbuf_size2_67_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_67_sram_inv[0:1]),
		.out(chanx_left_out_67_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_69 (
		.in({left_top_grid_pin_37_[0], chany_top_in_53_[0]}),
		.sram(mux_tree_like_tapbuf_size2_68_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_68_sram_inv[0:1]),
		.out(chanx_left_out_69_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_71 (
		.in({left_top_grid_pin_38_[0], chany_top_in_51_[0]}),
		.sram(mux_tree_like_tapbuf_size2_69_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_69_sram_inv[0:1]),
		.out(chanx_left_out_71_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_73 (
		.in({left_top_grid_pin_39_[0], chany_top_in_49_[0]}),
		.sram(mux_tree_like_tapbuf_size2_70_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_70_sram_inv[0:1]),
		.out(chanx_left_out_73_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_75 (
		.in({left_bottom_grid_pin_1_[0], chany_top_in_47_[0]}),
		.sram(mux_tree_like_tapbuf_size2_71_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_71_sram_inv[0:1]),
		.out(chanx_left_out_75_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_81 (
		.in({left_top_grid_pin_35_[0], chany_top_in_41_[0]}),
		.sram(mux_tree_like_tapbuf_size2_72_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_72_sram_inv[0:1]),
		.out(chanx_left_out_81_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_83 (
		.in({left_top_grid_pin_36_[0], chany_top_in_39_[0]}),
		.sram(mux_tree_like_tapbuf_size2_73_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_73_sram_inv[0:1]),
		.out(chanx_left_out_83_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_85 (
		.in({left_top_grid_pin_37_[0], chany_top_in_37_[0]}),
		.sram(mux_tree_like_tapbuf_size2_74_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_74_sram_inv[0:1]),
		.out(chanx_left_out_85_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_87 (
		.in({left_top_grid_pin_38_[0], chany_top_in_35_[0]}),
		.sram(mux_tree_like_tapbuf_size2_75_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_75_sram_inv[0:1]),
		.out(chanx_left_out_87_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_89 (
		.in({left_top_grid_pin_39_[0], chany_top_in_33_[0]}),
		.sram(mux_tree_like_tapbuf_size2_76_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_76_sram_inv[0:1]),
		.out(chanx_left_out_89_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_91 (
		.in({left_bottom_grid_pin_1_[0], chany_top_in_31_[0]}),
		.sram(mux_tree_like_tapbuf_size2_77_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_77_sram_inv[0:1]),
		.out(chanx_left_out_91_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_97 (
		.in({left_top_grid_pin_35_[0], chany_top_in_25_[0]}),
		.sram(mux_tree_like_tapbuf_size2_78_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_78_sram_inv[0:1]),
		.out(chanx_left_out_97_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_99 (
		.in({left_top_grid_pin_36_[0], chany_top_in_23_[0]}),
		.sram(mux_tree_like_tapbuf_size2_79_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_79_sram_inv[0:1]),
		.out(chanx_left_out_99_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_101 (
		.in({left_top_grid_pin_37_[0], chany_top_in_21_[0]}),
		.sram(mux_tree_like_tapbuf_size2_80_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_80_sram_inv[0:1]),
		.out(chanx_left_out_101_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_103 (
		.in({left_top_grid_pin_38_[0], chany_top_in_19_[0]}),
		.sram(mux_tree_like_tapbuf_size2_81_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_81_sram_inv[0:1]),
		.out(chanx_left_out_103_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_105 (
		.in({left_top_grid_pin_39_[0], chany_top_in_17_[0]}),
		.sram(mux_tree_like_tapbuf_size2_82_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_82_sram_inv[0:1]),
		.out(chanx_left_out_105_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_107 (
		.in({left_bottom_grid_pin_1_[0], chany_top_in_15_[0]}),
		.sram(mux_tree_like_tapbuf_size2_83_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_83_sram_inv[0:1]),
		.out(chanx_left_out_107_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_113 (
		.in({left_top_grid_pin_35_[0], chany_top_in_9_[0]}),
		.sram(mux_tree_like_tapbuf_size2_84_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_84_sram_inv[0:1]),
		.out(chanx_left_out_113_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_115 (
		.in({left_top_grid_pin_36_[0], chany_top_in_7_[0]}),
		.sram(mux_tree_like_tapbuf_size2_85_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_85_sram_inv[0:1]),
		.out(chanx_left_out_115_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_117 (
		.in({left_top_grid_pin_37_[0], chany_top_in_5_[0]}),
		.sram(mux_tree_like_tapbuf_size2_86_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_86_sram_inv[0:1]),
		.out(chanx_left_out_117_[0]));

	mux_tree_like_tapbuf_size2 mux_left_track_119 (
		.in({left_top_grid_pin_38_[0], chany_top_in_3_[0]}),
		.sram(mux_tree_like_tapbuf_size2_87_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size2_87_sram_inv[0:1]),
		.out(chanx_left_out_119_[0]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_0 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(ccff_head[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_0_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_0_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_2 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_0_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_1_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_1_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_4 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_1_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_2_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_2_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_6 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_2_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_3_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_3_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_8 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_3_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_4_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_4_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_10 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_4_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_5_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_5_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_20 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size3_mem_1_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_6_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_6_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_22 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_6_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_7_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_7_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_24 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_7_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_8_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_8_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_26 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_8_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_9_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_9_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_32 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_9_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_10_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_10_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_34 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_10_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_11_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_11_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_36 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_11_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_12_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_12_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_38 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_12_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_13_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_13_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_40 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_13_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_14_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_14_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_42 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_14_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_15_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_15_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_48 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_15_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_16_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_16_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_16_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_50 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_16_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_17_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_17_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_17_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_52 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_17_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_18_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_18_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_18_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_54 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_18_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_19_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_19_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_19_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_56 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_19_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_20_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_20_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_20_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_58 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_20_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_21_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_21_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_21_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_64 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_21_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_22_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_22_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_22_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_66 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_22_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_23_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_23_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_23_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_68 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_23_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_24_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_24_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_24_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_70 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_24_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_25_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_25_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_25_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_72 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_25_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_26_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_26_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_26_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_74 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_26_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_27_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_27_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_27_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_80 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_27_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_28_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_28_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_28_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_82 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_28_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_29_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_29_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_29_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_84 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_29_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_30_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_30_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_30_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_86 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_30_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_31_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_31_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_31_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_88 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_31_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_32_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_32_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_32_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_90 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_32_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_33_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_33_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_33_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_96 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_33_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_34_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_34_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_34_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_98 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_34_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_35_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_35_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_35_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_100 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_35_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_36_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_36_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_36_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_102 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_36_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_37_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_37_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_37_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_104 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_37_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_38_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_38_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_38_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_106 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_38_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_39_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_39_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_39_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_112 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_39_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_40_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_40_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_40_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_114 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_40_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_41_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_41_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_41_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_116 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_41_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_42_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_42_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_42_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_top_track_118 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_42_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_43_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_43_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_43_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_1 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_43_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_44_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_44_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_44_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_3 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_44_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_45_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_45_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_45_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_5 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_45_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_46_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_46_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_46_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_7 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_46_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_47_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_47_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_47_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_9 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_47_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_48_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_48_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_48_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_11 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_48_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_49_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_49_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_49_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_21 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size3_mem_3_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_50_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_50_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_50_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_23 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_50_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_51_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_51_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_51_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_25 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_51_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_52_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_52_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_52_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_27 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_52_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_53_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_53_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_53_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_33 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_53_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_54_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_54_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_54_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_35 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_54_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_55_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_55_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_55_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_37 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_55_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_56_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_56_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_56_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_39 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_56_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_57_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_57_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_57_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_41 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_57_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_58_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_58_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_58_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_43 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_58_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_59_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_59_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_59_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_49 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_59_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_60_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_60_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_60_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_51 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_60_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_61_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_61_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_61_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_53 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_61_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_62_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_62_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_62_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_55 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_62_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_63_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_63_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_63_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_57 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_63_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_64_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_64_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_64_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_59 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_64_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_65_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_65_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_65_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_65 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_65_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_66_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_66_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_66_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_67 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_66_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_67_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_67_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_67_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_69 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_67_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_68_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_68_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_68_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_71 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_68_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_69_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_69_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_69_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_73 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_69_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_70_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_70_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_70_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_75 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_70_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_71_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_71_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_71_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_81 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_71_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_72_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_72_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_72_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_83 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_72_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_73_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_73_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_73_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_85 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_73_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_74_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_74_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_74_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_87 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_74_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_75_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_75_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_75_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_89 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_75_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_76_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_76_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_76_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_91 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_76_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_77_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_77_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_77_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_97 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_77_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_78_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_78_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_78_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_99 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_78_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_79_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_79_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_79_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_101 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_79_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_80_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_80_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_80_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_103 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_80_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_81_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_81_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_81_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_105 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_81_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_82_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_82_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_82_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_107 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_82_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_83_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_83_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_83_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_113 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_83_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_84_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_84_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_84_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_115 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_84_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_85_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_85_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_85_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_117 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_85_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size2_mem_86_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_86_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_86_sram_inv[0:1]));

	mux_tree_like_tapbuf_size2_mem mem_left_track_119 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_86_ccff_tail[0]),
		.ccff_tail(ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size2_87_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size2_87_sram_inv[0:1]));

	mux_tree_like_tapbuf_size3 mux_top_track_16 (
		.in({top_left_grid_pin_30_[0], top_left_grid_pin_34_[0], chanx_left_in_104_[0]}),
		.sram(mux_tree_like_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size3_0_sram_inv[0:1]),
		.out(chany_top_out_16_[0]));

	mux_tree_like_tapbuf_size3 mux_top_track_18 (
		.in({top_left_grid_pin_31_[0], top_right_grid_pin_1_[0], chanx_left_in_102_[0]}),
		.sram(mux_tree_like_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size3_1_sram_inv[0:1]),
		.out(chany_top_out_18_[0]));

	mux_tree_like_tapbuf_size3 mux_left_track_17 (
		.in({left_top_grid_pin_35_[0], left_top_grid_pin_39_[0], chany_top_in_105_[0]}),
		.sram(mux_tree_like_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size3_2_sram_inv[0:1]),
		.out(chanx_left_out_17_[0]));

	mux_tree_like_tapbuf_size3 mux_left_track_19 (
		.in({left_top_grid_pin_36_[0], left_bottom_grid_pin_1_[0], chany_top_in_103_[0]}),
		.sram(mux_tree_like_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_tree_like_tapbuf_size3_3_sram_inv[0:1]),
		.out(chanx_left_out_19_[0]));

	mux_tree_like_tapbuf_size3_mem mem_top_track_16 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_5_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size3_mem_0_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size3_0_sram_inv[0:1]));

	mux_tree_like_tapbuf_size3_mem mem_top_track_18 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size3_mem_0_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size3_mem_1_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size3_1_sram_inv[0:1]));

	mux_tree_like_tapbuf_size3_mem mem_left_track_17 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size2_mem_49_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size3_mem_2_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size3_2_sram_inv[0:1]));

	mux_tree_like_tapbuf_size3_mem mem_left_track_19 (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.ccff_head(mux_tree_like_tapbuf_size3_mem_2_ccff_tail[0]),
		.ccff_tail(mux_tree_like_tapbuf_size3_mem_3_ccff_tail[0]),
		.mem_out(mux_tree_like_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_tree_like_tapbuf_size3_3_sram_inv[0:1]));

endmodule
// ----- END Verilog module for sb_22__0_ -----


