magic
tech sky130A
magscale 1 2
timestamp 1636140361
<< checkpaint >>
rect 39894 53320 48514 57324
<< locali >>
rect 47204 56044 47238 56060
rect 47204 55994 47238 56010
rect 47204 54634 47238 54650
rect 47204 54584 47238 54600
<< viali >>
rect 47204 56010 47238 56044
rect 47204 54600 47238 54634
<< metal1 >>
rect 47189 56001 47195 56053
rect 47247 56001 47253 56053
rect 47189 54591 47195 54643
rect 47247 54591 47253 54643
<< via1 >>
rect 47195 56044 47247 56053
rect 47195 56010 47204 56044
rect 47204 56010 47238 56044
rect 47238 56010 47247 56044
rect 47195 56001 47247 56010
rect 47195 54634 47247 54643
rect 47195 54600 47204 54634
rect 47204 54600 47238 54634
rect 47238 54600 47247 54634
rect 47195 54591 47247 54600
<< metal2 >>
rect 46666 56055 46722 56064
rect 46666 55990 46722 55999
rect 47193 56055 47249 56064
rect 47193 55990 47249 55999
rect 46680 55017 46708 55990
rect 46666 55008 46722 55017
rect 46666 54943 46722 54952
rect 46802 54884 46858 54893
rect 46802 54819 46858 54828
rect 46816 54654 46844 54819
rect 46802 54645 46858 54654
rect 46802 54580 46858 54589
rect 47193 54645 47249 54654
rect 47193 54580 47249 54589
<< via2 >>
rect 46666 55999 46722 56055
rect 47193 56053 47249 56055
rect 47193 56001 47195 56053
rect 47195 56001 47247 56053
rect 47247 56001 47249 56053
rect 47193 55999 47249 56001
rect 46666 54952 46722 55008
rect 46802 54828 46858 54884
rect 46802 54589 46858 54645
rect 47193 54643 47249 54645
rect 47193 54591 47195 54643
rect 47195 54591 47247 54643
rect 47247 54591 47249 54643
rect 47193 54589 47249 54591
<< metal3 >>
rect 46661 56057 46727 56060
rect 47188 56057 47254 56060
rect 46661 56055 47254 56057
rect 46661 55999 46666 56055
rect 46722 55999 47193 56055
rect 47249 55999 47254 56055
rect 46661 55997 47254 55999
rect 46661 55994 46727 55997
rect 47188 55994 47254 55997
rect 46661 55010 46727 55013
rect 41154 55008 46727 55010
rect 41154 54952 46666 55008
rect 46722 54952 46727 55008
rect 41154 54950 46727 54952
rect 46661 54947 46727 54950
rect 46797 54886 46863 54889
rect 41154 54884 46863 54886
rect 41154 54828 46802 54884
rect 46858 54828 46863 54884
rect 41154 54826 46863 54828
rect 46797 54823 46863 54826
rect 46797 54647 46863 54650
rect 47188 54647 47254 54650
rect 46797 54645 47254 54647
rect 46797 54589 46802 54645
rect 46858 54589 47193 54645
rect 47249 54589 47254 54645
rect 46797 54587 47254 54589
rect 46797 54584 46863 54587
rect 47188 54584 47254 54587
use contact_9  contact_9_0
timestamp 1636140361
transform 1 0 46797 0 1 54819
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1636140361
transform 1 0 47188 0 1 54580
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1636140361
transform 1 0 47189 0 1 54585
box 0 0 1 1
use contact_7  contact_7_0
timestamp 1636140361
transform 1 0 47192 0 1 54584
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1636140361
transform 1 0 46797 0 1 54580
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1636140361
transform 1 0 46661 0 1 54943
box 0 0 1 1
use contact_9  contact_9_4
timestamp 1636140361
transform 1 0 47188 0 1 55990
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1636140361
transform 1 0 47189 0 1 55995
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1636140361
transform 1 0 47192 0 1 55994
box 0 0 1 1
use contact_9  contact_9_5
timestamp 1636140361
transform 1 0 46661 0 1 55990
box 0 0 1 1
<< properties >>
string FIXED_BBOX 41154 54580 47254 56064
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_END 4737612
string GDS_START 4736372
<< end >>
