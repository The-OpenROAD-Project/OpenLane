VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO efs8hd_a2111oi_2
   CLASS CORE ;
   FOREIGN efs8hd_a2111oi_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.5200 BY 3.4000 ;
   SITE unitehd ;
   PIN D1
      PORT
         LAYER li1 ;
	    RECT 0.6050 1.3450 1.4250 1.6150 ;
      END
   END D1
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 1.9850 1.1050 2.8550 1.6150 ;
      END
   END B1
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 3.8250 1.1050 4.7250 1.6150 ;
      END
   END A2
   PIN C1
      PORT
         LAYER li1 ;
	    RECT 0.1250 1.7850 1.8000 2.1000 ;
	    RECT 0.1250 1.3050 0.4350 1.7850 ;
	    RECT 1.6150 1.6200 1.8000 1.7850 ;
	    RECT 1.6150 1.2900 1.8150 1.6200 ;
      END
   END C1
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.9000 2.3150 2.1400 2.6300 ;
	    RECT 1.9700 2.0300 2.1400 2.3150 ;
	    RECT 1.9700 1.8050 3.2550 2.0300 ;
	    RECT 3.0250 0.9350 3.2550 1.8050 ;
	    RECT 0.0950 0.7650 5.3550 0.9350 ;
	    RECT 0.0950 0.3200 0.3800 0.7650 ;
	    RECT 1.0150 0.3200 1.2950 0.7650 ;
	    RECT 1.9650 0.3200 2.2950 0.7650 ;
	    RECT 2.9650 0.3450 3.2950 0.7650 ;
	    RECT 5.0200 0.3700 5.3550 0.7650 ;
      END
   END Y
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 3.4650 1.7850 5.2900 2.0950 ;
	    RECT 3.4650 1.2300 3.6550 1.7850 ;
	    RECT 4.8950 1.2450 5.2900 1.7850 ;
      END
   END A1
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5500 0.1050 0.8450 0.5950 ;
	    RECT 1.4650 0.1050 1.7950 0.5550 ;
	    RECT 2.4650 0.1050 2.7950 0.5550 ;
	    RECT 4.1250 0.1050 4.4550 0.5550 ;
	    RECT 0.5500 0.0850 4.4550 0.1050 ;
	    RECT 0.0000 -0.0850 5.5200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.5200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.5200 3.4850 ;
	    RECT 3.6900 3.2950 4.9000 3.3150 ;
	    RECT 3.6900 2.8450 4.0200 3.2950 ;
	    RECT 4.5700 2.8450 4.9000 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.5200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0950 2.8700 2.9850 3.0800 ;
	    RECT 0.0950 2.8450 2.1850 2.8700 ;
	    RECT 0.0950 2.3400 0.4600 2.8450 ;
	    RECT 2.8150 2.6700 2.9850 2.8700 ;
	    RECT 3.1550 2.6200 3.5200 3.0800 ;
	    RECT 4.1900 2.6300 4.4000 3.0800 ;
	    RECT 5.0700 2.6300 5.4000 3.0800 ;
	    RECT 4.1900 2.6200 5.4000 2.6300 ;
	    RECT 2.3100 2.4550 2.6400 2.5750 ;
	    RECT 3.1550 2.4550 5.4000 2.6200 ;
	    RECT 2.3100 2.3050 5.4000 2.4550 ;
	    RECT 2.3100 2.2450 3.3350 2.3050 ;
   END
END efs8hd_a2111oi_2

MACRO efs8hd_a211oi_2
   CLASS CORE ;
   FOREIGN efs8hd_a211oi_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.6000 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5750 2.2300 0.9050 2.6300 ;
	    RECT 0.5750 0.9350 0.8550 2.2300 ;
	    RECT 0.5750 0.7650 3.1450 0.9350 ;
	    RECT 0.5750 0.3200 0.8350 0.7650 ;
	    RECT 1.5050 0.3550 1.6950 0.7650 ;
      END
   END Y
   PIN C1
      PORT
         LAYER li1 ;
	    RECT 0.1000 1.1050 0.4050 2.0200 ;
      END
   END C1
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 1.0350 1.6150 1.2550 2.0200 ;
	    RECT 1.0350 1.2950 1.7850 1.6150 ;
      END
   END B1
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 2.3700 1.1050 3.0800 1.6150 ;
      END
   END A1
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 4.1750 1.6150 4.5000 2.0700 ;
	    RECT 3.7400 1.2950 4.5000 1.6150 ;
      END
   END A2
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1450 0.1050 0.3950 0.9350 ;
	    RECT 1.0050 0.1050 1.3350 0.5950 ;
	    RECT 1.8650 0.1050 2.1950 0.5950 ;
	    RECT 3.6750 0.1050 4.0050 0.5700 ;
	    RECT 0.1450 0.0850 4.0050 0.1050 ;
	    RECT 0.0000 -0.0850 4.6000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.6000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.6000 3.4850 ;
	    RECT 2.4350 3.2950 4.3850 3.3150 ;
	    RECT 2.4350 2.2950 2.6650 3.2950 ;
	    RECT 3.2950 2.2950 3.5250 3.2950 ;
	    RECT 4.1550 2.2950 4.3850 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.6000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1450 2.8550 2.2150 3.0700 ;
	    RECT 0.1450 2.2300 0.4050 2.8550 ;
	    RECT 1.0750 2.8200 2.2150 2.8550 ;
	    RECT 1.0750 2.2300 1.2650 2.8200 ;
	    RECT 1.4350 2.0700 1.7650 2.5950 ;
	    RECT 1.9350 2.2950 2.2150 2.8200 ;
	    RECT 2.8450 2.0700 3.1150 3.0800 ;
	    RECT 3.7050 2.0700 3.9750 3.0800 ;
	    RECT 1.4350 1.8200 3.9750 2.0700 ;
	    RECT 3.3250 0.7950 4.4350 1.0700 ;
	    RECT 3.3250 0.5950 3.4950 0.7950 ;
	    RECT 2.3850 0.3300 3.4950 0.5950 ;
	    RECT 4.1850 0.3300 4.4350 0.7950 ;
   END
END efs8hd_a211oi_2
MACRO efs8hd_a21boi_2
   CLASS CORE ;
   FOREIGN efs8hd_a21boi_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.1400 BY 3.4000 ;
   SITE unitehd ;
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 4.1400 3.5050 ;
	    RECT 0.0950 2.6000 0.4250 3.2950 ;
	    RECT 2.3850 2.7450 2.5550 3.2950 ;
	    RECT 3.1600 2.8450 3.4900 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.1400 3.7000 ;
      END
   END vpwr
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.9850 0.1050 1.2250 1.1050 ;
	    RECT 1.9400 0.1050 2.2700 0.5550 ;
	    RECT 3.6350 0.1050 3.9300 1.0800 ;
	    RECT 0.0000 -0.1050 4.1400 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.1400 0.3000 ;
      END
   END vgnd
   PIN B1N
      PORT
         LAYER li1 ;
	    RECT 0.1200 0.9550 0.4250 2.2550 ;
      END
   END B1N
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 2.1000 1.8700 3.6750 2.0950 ;
	    RECT 2.1000 1.5550 2.4250 1.8700 ;
	    RECT 2.0950 1.3450 2.4250 1.5550 ;
	    RECT 3.3850 1.6200 3.6750 1.8700 ;
	    RECT 3.3850 1.2950 3.7950 1.6200 ;
      END
   END A2
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 2.6050 1.2450 3.2150 1.6550 ;
      END
   END A1
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 1.5200 0.9800 1.7150 2.6450 ;
	    RECT 1.5200 0.7700 3.0600 0.9800 ;
	    RECT 1.5200 0.3200 1.7200 0.7700 ;
	    RECT 2.7300 0.3200 3.0600 0.7700 ;
      END
   END Y
   OBS
         LAYER li1 ;
	    RECT 1.0450 2.8550 2.2150 3.0800 ;
	    RECT 0.5950 1.6050 0.8550 2.8300 ;
	    RECT 1.0450 2.2450 1.3500 2.8550 ;
	    RECT 1.8850 2.5300 2.2150 2.8550 ;
	    RECT 2.8100 2.6300 2.9800 3.0800 ;
	    RECT 3.6600 2.6300 3.9200 3.0800 ;
	    RECT 2.8100 2.5300 3.9200 2.6300 ;
	    RECT 1.8850 2.3200 3.9200 2.5300 ;
	    RECT 0.5950 1.3400 1.3250 1.6050 ;
	    RECT 0.5950 0.6650 0.7950 1.3400 ;
	    RECT 0.2650 0.4500 0.7950 0.6650 ;
   END
END efs8hd_a21boi_2
MACRO efs8hd_a21oi_2
   CLASS CORE ;
   FOREIGN efs8hd_a21oi_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.2200 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 2.3150 0.9350 2.6150 2.6450 ;
	    RECT 0.9550 0.7650 2.6150 0.9350 ;
	    RECT 0.9550 0.3200 1.3000 0.7650 ;
	    RECT 2.2950 0.3200 2.6150 0.7650 ;
      END
   END Y
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 0.8150 1.1050 1.4250 1.6150 ;
      END
   END A1
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 2.8000 1.1050 3.0750 2.0300 ;
      END
   END B1
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 0.1450 1.7850 1.9300 2.0950 ;
	    RECT 0.1450 1.2950 0.6450 1.7850 ;
	    RECT 1.6050 1.5550 1.9300 1.7850 ;
	    RECT 1.6050 1.3450 1.9350 1.5550 ;
      END
   END A2
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1000 0.1050 0.3950 1.0800 ;
	    RECT 1.7600 0.1050 2.0900 0.5550 ;
	    RECT 2.7950 0.1050 3.1250 0.9350 ;
	    RECT 0.1000 0.0850 3.1250 0.1050 ;
	    RECT 0.0000 -0.0850 3.2200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.2200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.2200 3.4850 ;
	    RECT 0.5400 3.2950 1.6450 3.3150 ;
	    RECT 0.5400 2.8450 0.8700 3.2950 ;
	    RECT 1.4750 2.7450 1.6450 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.2200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1100 2.6300 0.3700 3.0800 ;
	    RECT 1.0500 2.6300 1.2200 3.0800 ;
	    RECT 0.1100 2.5300 1.2200 2.6300 ;
	    RECT 1.8150 2.8550 3.0900 3.0800 ;
	    RECT 1.8150 2.5300 2.1450 2.8550 ;
	    RECT 0.1100 2.3200 2.1450 2.5300 ;
	    RECT 2.7850 2.2450 3.0900 2.8550 ;
   END
END efs8hd_a21oi_2
MACRO efs8hd_a221oi_2
   CLASS CORE ;
   FOREIGN efs8hd_a221oi_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.5200 BY 3.4000 ;
   SITE unitehd ;
   PIN C1
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.3450 0.4200 2.0200 ;
      END
   END C1
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5950 1.1300 0.8450 2.6550 ;
	    RECT 0.5950 1.0800 4.3950 1.1300 ;
	    RECT 0.5150 0.9050 4.3950 1.0800 ;
	    RECT 0.5150 0.3800 0.8550 0.9050 ;
	    RECT 2.2850 0.8050 2.6350 0.9050 ;
	    RECT 4.0650 0.8050 4.3950 0.9050 ;
      END
   END Y
   PIN B2
      PORT
         LAYER li1 ;
	    RECT 1.5050 1.7850 3.2650 2.0200 ;
	    RECT 1.5050 1.3450 2.0400 1.7850 ;
	    RECT 2.9250 1.3450 3.2650 1.7850 ;
      END
   END B2
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 2.2100 1.3450 2.7550 1.6150 ;
      END
   END B1
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 3.8250 1.3450 4.4800 1.6150 ;
      END
   END A1
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 3.4350 1.7850 4.8200 2.0200 ;
	    RECT 3.4350 1.3050 3.6550 1.7850 ;
	    RECT 4.6500 1.6150 4.8200 1.7850 ;
	    RECT 4.6500 1.3450 5.4350 1.6150 ;
      END
   END A2
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1050 0.1050 0.3450 1.1200 ;
	    RECT 1.0250 0.1050 1.7050 0.6950 ;
	    RECT 3.2700 0.1050 3.4400 0.6950 ;
	    RECT 4.9850 0.1050 5.1550 1.1300 ;
	    RECT 0.1050 0.0850 5.1550 0.1050 ;
	    RECT 0.0000 -0.0850 5.5200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.5200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.5200 3.4850 ;
	    RECT 3.6850 3.2950 4.7750 3.3150 ;
	    RECT 3.6850 2.6550 3.9350 3.2950 ;
	    RECT 4.5250 2.6550 4.7750 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.5200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0900 2.8700 1.2750 3.0800 ;
	    RECT 0.0900 2.2450 0.4250 2.8700 ;
	    RECT 1.0150 2.4450 1.2750 2.8700 ;
	    RECT 1.5050 2.8700 3.4750 3.0800 ;
	    RECT 1.5050 2.6550 1.7550 2.8700 ;
	    RECT 2.3450 2.6550 2.5950 2.8700 ;
	    RECT 1.9250 2.4450 2.1750 2.6550 ;
	    RECT 2.7650 2.4450 3.0150 2.6550 ;
	    RECT 1.0150 2.2300 3.0150 2.4450 ;
	    RECT 3.2250 2.4450 3.4750 2.8700 ;
	    RECT 4.1050 2.4450 4.3550 3.0800 ;
	    RECT 4.9900 2.4450 5.1950 3.0800 ;
	    RECT 3.2250 2.2300 5.1950 2.4450 ;
	    RECT 1.0150 1.8700 1.2750 2.2300 ;
	    RECT 4.9900 1.8200 5.1950 2.2300 ;
	    RECT 4.5650 0.5950 4.8150 1.1300 ;
	    RECT 1.8750 0.3200 3.0550 0.5950 ;
	    RECT 3.6450 0.3200 4.8150 0.5950 ;
   END
END efs8hd_a221oi_2
MACRO efs8hd_a22oi_2
   CLASS CORE ;
   FOREIGN efs8hd_a22oi_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.6000 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.6400 ;
	    RECT 3.5550 0.1050 3.8850 0.6400 ;
	    RECT 0.5150 0.0850 3.8850 0.1050 ;
	    RECT 0.0000 -0.0850 4.6000 0.0850 ;
	    RECT 0.6100 -0.1050 0.7800 -0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.6000 0.3000 ;
      END
   END vgnd
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.0950 2.0700 0.3450 3.0800 ;
	    RECT 0.9350 2.0700 1.2650 2.6550 ;
	    RECT 1.7750 2.0700 2.1600 2.6550 ;
	    RECT 0.0950 1.8550 2.1600 2.0700 ;
	    RECT 1.8700 1.0550 2.1600 1.8550 ;
	    RECT 1.3550 0.8450 3.0450 1.0550 ;
      END
   END Y
   PIN B2
      PORT
         LAYER li1 ;
	    RECT 0.1450 1.3450 0.7800 1.6150 ;
      END
   END B2
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 1.0650 1.3450 1.7000 1.6150 ;
      END
   END B1
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 2.4450 1.3450 3.1000 1.6150 ;
      END
   END A1
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 3.3650 1.3450 4.5000 1.6150 ;
      END
   END A2
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.6100 3.4850 0.7800 3.5050 ;
	    RECT 0.0000 3.3150 4.6000 3.4850 ;
	    RECT 0.6100 3.2950 0.7800 3.3150 ;
	    RECT 2.7950 3.2950 3.8050 3.3150 ;
	    RECT 2.7950 2.2800 2.9650 3.2950 ;
	    RECT 3.6350 2.2800 3.8050 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.6000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.5150 2.8700 2.6250 3.0800 ;
	    RECT 0.5150 2.2800 0.7650 2.8700 ;
	    RECT 1.4350 2.2800 1.6050 2.8700 ;
	    RECT 2.3750 2.0700 2.6250 2.8700 ;
	    RECT 3.1350 2.0700 3.4650 3.0800 ;
	    RECT 3.9750 2.0700 4.3050 3.0800 ;
	    RECT 2.3750 1.8550 4.3050 2.0700 ;
	    RECT 0.0950 0.8500 1.1850 1.0650 ;
	    RECT 0.0950 0.3200 0.3450 0.8500 ;
	    RECT 1.0150 0.6300 1.1850 0.8500 ;
	    RECT 3.2150 0.8500 4.3750 1.0650 ;
	    RECT 3.2150 0.6300 3.3850 0.8500 ;
	    RECT 1.0150 0.3200 2.1050 0.6300 ;
	    RECT 2.2950 0.3200 3.3850 0.6300 ;
	    RECT 4.0550 0.3200 4.3750 0.8500 ;
   END
END efs8hd_a22oi_2
MACRO efs8hd_a2bb2oi_2
   CLASS CORE ;
   FOREIGN efs8hd_a2bb2oi_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.5200 BY 3.4000 ;
   SITE unitehd ;
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.7850 2.0300 2.0200 ;
	    RECT 0.0850 1.3450 0.7100 1.7850 ;
	    RECT 1.7000 1.3450 2.0300 1.7850 ;
      END
   END B1
   PIN B2
      PORT
         LAYER li1 ;
	    RECT 0.9400 1.3450 1.4800 1.6150 ;
      END
   END B2
   PIN A1N
      PORT
         LAYER li1 ;
	    RECT 3.3100 1.3450 4.1150 1.6150 ;
      END
   END A1N
   PIN A2N
      PORT
         LAYER li1 ;
	    RECT 4.2850 1.3450 5.4350 1.6150 ;
      END
   END A2N
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 2.3700 2.0750 2.6200 2.6550 ;
	    RECT 2.3700 1.1300 2.6600 2.0750 ;
	    RECT 1.0700 0.9050 2.6600 1.1300 ;
	    RECT 1.0700 0.8050 1.4000 0.9050 ;
	    RECT 2.3300 0.3200 2.6600 0.9050 ;
      END
   END Y
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.3100 0.1050 0.4800 1.1200 ;
	    RECT 1.9900 0.1050 2.1600 0.6950 ;
	    RECT 2.8300 0.1050 3.5200 0.6950 ;
	    RECT 4.1900 0.1050 4.3600 0.6950 ;
	    RECT 5.0300 0.1050 5.2000 1.1300 ;
	    RECT 0.3100 0.0850 5.2000 0.1050 ;
	    RECT 0.0000 -0.0850 5.5200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.5200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.5200 3.4850 ;
	    RECT 0.6900 3.2950 3.9800 3.3150 ;
	    RECT 0.6900 2.6700 0.9400 3.2950 ;
	    RECT 1.5300 2.6700 1.7800 3.2950 ;
	    RECT 3.7300 2.6700 3.9800 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.5200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.2700 2.4450 0.5200 3.0800 ;
	    RECT 1.1100 2.4450 1.3600 3.0800 ;
	    RECT 1.9500 2.8700 3.0400 3.0800 ;
	    RECT 1.9500 2.4450 2.2000 2.8700 ;
	    RECT 0.2700 2.2300 2.2000 2.4450 ;
	    RECT 2.7900 2.2450 3.0400 2.8700 ;
	    RECT 3.3100 2.4550 3.5600 3.0800 ;
	    RECT 4.1500 2.8700 5.2400 3.0800 ;
	    RECT 4.1500 2.4550 4.4000 2.8700 ;
	    RECT 3.3100 2.2300 4.4000 2.4550 ;
	    RECT 4.5700 2.0200 4.8200 2.6550 ;
	    RECT 2.9500 1.8050 4.8200 2.0200 ;
	    RECT 4.9900 1.8200 5.2400 2.8700 ;
	    RECT 2.9500 1.6550 3.1200 1.8050 ;
	    RECT 2.8300 1.2450 3.1200 1.6550 ;
	    RECT 2.9500 1.1300 3.1200 1.2450 ;
	    RECT 0.6500 0.5950 0.9000 1.1200 ;
	    RECT 2.9500 0.9050 4.8600 1.1300 ;
	    RECT 0.6500 0.3200 1.8200 0.5950 ;
	    RECT 3.6900 0.3200 4.0200 0.9050 ;
	    RECT 4.5300 0.3200 4.8600 0.9050 ;
   END
END efs8hd_a2bb2oi_2
MACRO efs8hd_a311oi_2
   CLASS CORE ;
   FOREIGN efs8hd_a311oi_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.5200 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 4.6600 2.3950 5.0050 2.6050 ;
	    RECT 4.6600 2.1800 4.9900 2.3950 ;
	    RECT 4.6600 2.1000 5.0050 2.1800 ;
	    RECT 4.2600 1.9700 5.0050 2.1000 ;
	    RECT 4.2600 1.8900 4.9900 1.9700 ;
	    RECT 4.2600 1.0300 4.4750 1.8900 ;
	    RECT 4.2600 0.9350 5.3450 1.0300 ;
	    RECT 2.2950 0.7650 5.3450 0.9350 ;
	    RECT 3.2350 0.3200 3.4050 0.7650 ;
	    RECT 4.0850 0.3200 4.2550 0.7650 ;
	    RECT 5.1750 0.3200 5.3450 0.7650 ;
      END
   END Y
   PIN A3
      PORT
         LAYER li1 ;
	    RECT 0.1350 1.1050 0.8000 1.6550 ;
      END
   END A3
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 1.0550 1.1050 1.8050 1.6550 ;
      END
   END A2
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 1.9850 1.2450 3.1150 1.6550 ;
      END
   END A1
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 3.3650 1.1050 4.0550 1.6550 ;
      END
   END B1
   PIN C1
      PORT
         LAYER li1 ;
	    RECT 5.1750 1.6200 5.4100 2.0300 ;
	    RECT 4.7300 1.3450 5.4100 1.6200 ;
      END
   END C1
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 3.5850 0.1050 3.9150 0.5800 ;
	    RECT 4.6750 0.1050 5.0050 0.5800 ;
	    RECT 0.5150 0.0850 5.0050 0.1050 ;
	    RECT 0.0000 -0.0850 5.5200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.5200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.5200 3.4850 ;
	    RECT 0.0950 3.2950 2.9750 3.3150 ;
	    RECT 0.0950 1.8700 0.3450 3.2950 ;
	    RECT 0.9350 2.3950 1.2650 3.2950 ;
	    RECT 1.7850 2.3950 2.1350 3.2950 ;
	    RECT 2.6450 2.3950 2.9750 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.5200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.5950 2.1800 0.7650 3.0800 ;
	    RECT 1.4350 2.1800 1.6050 3.0800 ;
	    RECT 2.3050 2.1800 2.4750 3.0800 ;
	    RECT 4.1100 3.0300 4.4400 3.0800 ;
	    RECT 5.1750 3.0300 5.3450 3.0800 ;
	    RECT 3.1450 2.8200 5.3450 3.0300 ;
	    RECT 3.5850 2.1800 3.9150 2.6050 ;
	    RECT 4.1100 2.3950 4.4400 2.8200 ;
	    RECT 5.1750 2.2450 5.3450 2.8200 ;
	    RECT 0.5950 1.9700 3.9150 2.1800 ;
	    RECT 0.1750 0.7650 2.1050 0.9350 ;
	    RECT 0.1750 0.3200 0.3450 0.7650 ;
	    RECT 1.0150 0.3200 1.1850 0.7650 ;
	    RECT 1.3550 0.3800 3.0450 0.5950 ;
   END
END efs8hd_a311oi_2
MACRO efs8hd_a31oi_2
   CLASS CORE ;
   FOREIGN efs8hd_a31oi_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.6000 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 3.7550 2.0200 4.0850 2.6450 ;
	    RECT 3.2550 1.8050 4.0850 2.0200 ;
	    RECT 3.2550 1.0300 3.5700 1.8050 ;
	    RECT 2.2950 0.8200 4.5050 1.0300 ;
	    RECT 3.2550 0.3200 3.4250 0.8200 ;
	    RECT 4.1750 0.3700 4.5050 0.8200 ;
      END
   END Y
   PIN A3
      PORT
         LAYER li1 ;
	    RECT 0.1450 1.2450 0.8200 2.0200 ;
      END
   END A3
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 1.0500 1.2450 1.7550 2.0200 ;
      END
   END A2
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 1.9550 1.2450 2.6650 2.0200 ;
	    RECT 2.9050 1.2450 3.0750 1.6550 ;
      END
   END A1
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 4.2650 1.6150 4.4900 2.0300 ;
	    RECT 3.8200 1.3450 4.4900 1.6150 ;
      END
   END B1
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 3.6750 0.1050 4.0050 0.5800 ;
	    RECT 0.5150 0.0850 4.0050 0.1050 ;
	    RECT 0.0000 -0.0850 4.6000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.6000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.6000 3.4850 ;
	    RECT 0.5150 3.2950 2.9800 3.3150 ;
	    RECT 0.5150 2.6550 0.8450 3.2950 ;
	    RECT 1.3550 2.6550 1.6850 3.2950 ;
	    RECT 2.3100 2.6550 2.9800 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.6000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1750 2.4450 0.3450 3.0800 ;
	    RECT 1.0150 2.4450 1.1850 3.0800 ;
	    RECT 1.8550 2.4450 2.0250 3.0800 ;
	    RECT 3.3350 2.8700 4.4250 3.0800 ;
	    RECT 3.3350 2.4450 3.5050 2.8700 ;
	    RECT 0.1750 2.2300 3.5050 2.4450 ;
	    RECT 4.2550 2.2450 4.4250 2.8700 ;
	    RECT 0.0950 0.8200 2.1050 1.0300 ;
	    RECT 1.3550 0.3700 3.0750 0.5800 ;
   END
END efs8hd_a31oi_2
MACRO efs8hd_and2_2
   CLASS CORE ;
   FOREIGN efs8hd_and2_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 2.7600 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 1.7650 2.3950 2.2150 3.0800 ;
	    RECT 1.9650 0.6800 2.2150 2.3950 ;
	    RECT 1.6650 0.3200 2.2150 0.6800 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.6550 0.4000 2.2050 ;
	    RECT 0.0850 1.3450 0.7750 1.6550 ;
      END
   END A
   PIN B
      PORT
         LAYER li1 ;
	    RECT 1.0050 1.3450 1.3350 1.6550 ;
      END
   END B
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 1.2450 0.1050 1.4950 0.6800 ;
	    RECT 2.3850 0.1050 2.6750 1.1050 ;
	    RECT 1.2450 0.0850 2.6750 0.1050 ;
	    RECT 0.0000 -0.0850 2.7600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 2.7600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 2.7600 3.4850 ;
	    RECT 0.2850 3.2950 2.6750 3.3150 ;
	    RECT 0.2850 2.4550 0.5650 3.2950 ;
	    RECT 1.2450 2.3950 1.5750 3.2950 ;
	    RECT 2.3850 1.8700 2.6750 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 2.7600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.7350 2.1800 1.0350 2.8700 ;
	    RECT 0.7350 1.9700 1.6750 2.1800 ;
	    RECT 1.5050 1.6550 1.6750 1.9700 ;
	    RECT 1.5050 1.2450 1.7950 1.6550 ;
	    RECT 1.5050 1.1300 1.6750 1.2450 ;
	    RECT 0.2850 0.8950 1.6750 1.1300 ;
	    RECT 0.2850 0.4450 0.6150 0.8950 ;
   END
END efs8hd_and2_2
MACRO efs8hd_and2b_2
   CLASS CORE ;
   FOREIGN efs8hd_and2b_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.2200 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 2.3750 1.9750 2.6800 2.9550 ;
	    RECT 2.5050 0.9700 2.6800 1.9750 ;
	    RECT 2.4450 0.3200 2.6800 0.9700 ;
      END
   END X
   PIN AN
      PORT
         LAYER li1 ;
	    RECT 0.1450 0.9550 0.4500 2.0200 ;
      END
   END AN
   PIN B
      PORT
         LAYER li1 ;
	    RECT 1.5050 2.0550 2.2000 2.6350 ;
      END
   END B
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0950 0.1050 0.4250 0.7400 ;
	    RECT 1.8750 0.1050 2.2750 0.7250 ;
	    RECT 2.8650 0.1050 3.1350 0.9000 ;
	    RECT 0.0950 0.0850 3.1350 0.1050 ;
	    RECT 0.0000 -0.0850 3.2200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.2200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.2200 3.4850 ;
	    RECT 0.5150 3.2950 3.1350 3.3150 ;
	    RECT 0.5150 2.7300 0.8450 3.2950 ;
	    RECT 1.5100 2.8050 2.1950 3.2950 ;
	    RECT 2.8650 2.1000 3.1350 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.2200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1750 2.5200 0.3450 3.0550 ;
	    RECT 0.1750 2.2300 0.8550 2.5200 ;
	    RECT 0.6200 1.4200 0.8550 2.2300 ;
	    RECT 1.0450 1.8450 1.3300 3.0250 ;
	    RECT 1.0450 1.6550 1.9050 1.8450 ;
	    RECT 1.0450 1.6300 2.3350 1.6550 ;
	    RECT 0.6200 1.0050 1.1750 1.4200 ;
	    RECT 1.3450 1.1800 2.3350 1.6300 ;
	    RECT 0.6200 0.8200 0.8350 1.0050 ;
	    RECT 0.5950 0.3500 0.8350 0.8200 ;
	    RECT 1.3450 0.7650 1.5150 1.1800 ;
	    RECT 1.1150 0.5200 1.5150 0.7650 ;
	    RECT 1.1150 0.3400 1.2850 0.5200 ;
   END
END efs8hd_and2b_2
MACRO efs8hd_and3_2
   CLASS CORE ;
   FOREIGN efs8hd_and3_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 2.7600 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 1.9700 2.2450 2.2450 3.0800 ;
	    RECT 2.0750 1.8050 2.2450 2.2450 ;
	    RECT 2.0600 1.1550 2.6750 1.8050 ;
	    RECT 2.0600 0.8950 2.2300 1.1550 ;
	    RECT 1.9800 0.3200 2.2300 0.8950 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.7650 0.4700 1.6150 ;
      END
   END A
   PIN C
      PORT
         LAYER li1 ;
	    RECT 1.0650 0.9400 1.4750 1.5550 ;
	    RECT 1.0650 0.3800 1.2950 0.9400 ;
      END
   END C
   PIN B
      PORT
         LAYER li1 ;
	    RECT 0.9450 2.4650 1.3700 3.0800 ;
      END
   END B
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 1.4750 0.1050 1.8050 0.7250 ;
	    RECT 2.4000 0.1050 2.6750 0.9300 ;
	    RECT 1.4750 0.0850 2.6750 0.1050 ;
	    RECT 0.0000 -0.0850 2.7600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 2.7600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 2.7600 3.4850 ;
	    RECT 0.0850 3.2950 2.6750 3.3150 ;
	    RECT 0.0850 2.6650 0.7150 3.2950 ;
	    RECT 0.5250 2.4950 0.7150 2.6650 ;
	    RECT 0.5250 2.1650 0.7750 2.4950 ;
	    RECT 1.5550 2.2400 1.7700 3.2950 ;
	    RECT 2.4150 2.0300 2.6750 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 2.7600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1000 1.9950 0.3550 2.4500 ;
	    RECT 1.0800 1.9950 1.3300 2.2950 ;
	    RECT 0.1000 1.7850 1.8900 1.9950 ;
	    RECT 0.6400 1.7800 1.8900 1.7850 ;
	    RECT 0.6400 0.5950 0.8950 1.7800 ;
	    RECT 1.6600 1.2450 1.8900 1.7800 ;
	    RECT 0.1050 0.3800 0.8950 0.5950 ;
   END
END efs8hd_and3_2
MACRO efs8hd_and3b_2
   CLASS CORE ;
   FOREIGN efs8hd_and3b_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.6800 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 2.8750 2.2450 3.1600 3.0800 ;
	    RECT 2.9900 1.8050 3.1600 2.2450 ;
	    RECT 2.9900 1.1550 3.5950 1.8050 ;
	    RECT 2.9900 0.8950 3.1600 1.1550 ;
	    RECT 2.9150 0.3200 3.1600 0.8950 ;
      END
   END X
   PIN C
      PORT
         LAYER li1 ;
	    RECT 1.9850 0.9550 2.4200 1.5550 ;
	    RECT 1.9850 0.3800 2.2200 0.9550 ;
      END
   END C
   PIN AN
      PORT
         LAYER li1 ;
	    RECT 0.1450 0.7650 0.4100 1.6550 ;
      END
   END AN
   PIN B
      PORT
         LAYER li1 ;
	    RECT 1.8150 2.4650 2.2900 3.0800 ;
      END
   END B
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.1050 0.4250 0.5950 ;
	    RECT 2.4100 0.1050 2.7400 0.7250 ;
	    RECT 3.3300 0.1050 3.5950 0.9300 ;
	    RECT 0.0850 0.0850 3.5950 0.1050 ;
	    RECT 0.0000 -0.0850 3.6800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.6800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.6800 3.4850 ;
	    RECT 0.0850 3.2950 3.5950 3.3150 ;
	    RECT 0.0850 1.9700 0.4000 3.2950 ;
	    RECT 1.0300 2.6650 1.6450 3.2950 ;
	    RECT 1.4550 2.2950 1.6450 2.6650 ;
	    RECT 1.4550 2.1250 1.7850 2.2950 ;
	    RECT 2.4600 2.2400 2.6750 3.2950 ;
	    RECT 3.3300 2.0300 3.5950 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.6800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.5950 1.5550 0.8550 2.3800 ;
	    RECT 1.0500 1.9550 1.2850 2.4500 ;
	    RECT 2.0100 1.9950 2.2000 2.2950 ;
	    RECT 2.0100 1.9550 2.8200 1.9950 ;
	    RECT 1.0500 1.7800 2.8200 1.9550 ;
	    RECT 0.5950 1.2700 1.4150 1.5550 ;
	    RECT 0.5950 0.3800 0.8550 1.2700 ;
	    RECT 1.5850 0.7150 1.8150 1.7800 ;
	    RECT 2.5900 1.2450 2.8200 1.7800 ;
	    RECT 1.0550 0.3800 1.8150 0.7150 ;
   END
END efs8hd_and3b_2
MACRO efs8hd_and4_2
   CLASS CORE ;
   FOREIGN efs8hd_and4_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.6800 BY 3.4000 ;
   SITE unitehd ;
   PIN B
      PORT
         LAYER li1 ;
	    RECT 0.8900 0.5250 1.2450 1.6550 ;
      END
   END B
   PIN C
      PORT
         LAYER li1 ;
	    RECT 1.4200 1.6300 1.5900 1.6550 ;
	    RECT 1.4200 0.5200 1.7200 1.6300 ;
      END
   END C
   PIN X
      PORT
         LAYER li1 ;
	    RECT 2.7350 1.8700 3.0750 3.0800 ;
	    RECT 2.8950 1.0050 3.0750 1.8700 ;
	    RECT 2.7350 0.4250 3.0750 1.0050 ;
	    RECT 2.7350 0.3700 3.0650 0.4250 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.1250 0.9450 0.3300 2.5950 ;
      END
   END A
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.9000 0.5200 2.1600 1.6550 ;
      END
   END D
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 2.3300 0.1050 2.5650 1.1150 ;
	    RECT 3.2550 0.1050 3.5850 1.0150 ;
	    RECT 2.3300 0.0850 3.5850 0.1050 ;
	    RECT 0.0000 -0.0850 3.6800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.6800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.6800 3.4850 ;
	    RECT 0.0950 3.2950 3.5750 3.3150 ;
	    RECT 0.0950 2.8200 0.4250 3.2950 ;
	    RECT 1.0700 2.3950 1.4000 3.2950 ;
	    RECT 2.2350 2.2950 2.5650 3.2950 ;
	    RECT 3.2450 2.2950 3.5750 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.6800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.6000 2.0800 0.8500 3.0800 ;
	    RECT 1.5850 2.0800 1.8350 3.0800 ;
	    RECT 0.5000 1.8700 2.5550 2.0800 ;
	    RECT 0.5000 0.7300 0.6700 1.8700 ;
	    RECT 2.3300 1.6450 2.5550 1.8700 ;
	    RECT 2.3300 1.3450 2.7250 1.6450 ;
	    RECT 0.1750 0.3200 0.6700 0.7300 ;
   END
END efs8hd_and4_2
MACRO efs8hd_and4b_2
   CLASS CORE ;
   FOREIGN efs8hd_and4b_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.1400 BY 3.4000 ;
   SITE unitehd ;
   PIN B
      PORT
         LAYER li1 ;
	    RECT 1.5250 0.5250 1.7450 2.1800 ;
      END
   END B
   PIN C
      PORT
         LAYER li1 ;
	    RECT 1.9600 0.5250 2.2750 2.1200 ;
      END
   END C
   PIN X
      PORT
         LAYER li1 ;
	    RECT 3.3400 2.1800 3.5450 3.0800 ;
	    RECT 3.3400 1.9200 4.0550 2.1800 ;
	    RECT 3.4250 1.0300 4.0550 1.9200 ;
	    RECT 3.2600 0.8000 4.0550 1.0300 ;
	    RECT 3.2600 0.3200 3.5450 0.8000 ;
      END
   END X
   PIN AN
      PORT
         LAYER li1 ;
	    RECT 0.1350 0.9250 0.3350 2.0400 ;
      END
   END AN
   PIN D
      PORT
         LAYER li1 ;
	    RECT 2.4450 0.8050 2.7750 2.0200 ;
      END
   END D
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0950 0.1050 0.4250 0.5800 ;
	    RECT 2.7600 0.1050 3.0900 0.5800 ;
	    RECT 3.7150 0.1050 4.0500 0.5800 ;
	    RECT 0.0950 0.0850 4.0500 0.1050 ;
	    RECT 0.0000 -0.0850 4.1400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.1400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.1400 3.4850 ;
	    RECT 0.5150 3.2950 4.0500 3.3150 ;
	    RECT 0.5150 2.7450 0.8450 3.2950 ;
	    RECT 1.5550 2.8200 2.2250 3.2950 ;
	    RECT 2.8400 2.7450 3.1700 3.2950 ;
	    RECT 3.7150 2.3950 4.0500 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.1400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1750 2.5000 0.3450 3.0800 ;
	    RECT 1.0150 2.6050 1.1850 3.0800 ;
	    RECT 2.4400 2.6050 2.6100 3.0800 ;
	    RECT 0.1750 2.2900 0.8050 2.5000 ;
	    RECT 0.6350 1.6550 0.8050 2.2900 ;
	    RECT 1.0150 2.4550 2.6100 2.6050 ;
	    RECT 1.0150 2.3950 3.1650 2.4550 ;
	    RECT 1.0150 2.0750 1.3150 2.3950 ;
	    RECT 2.4400 2.2450 3.1650 2.3950 ;
	    RECT 0.6350 1.2450 0.9750 1.6550 ;
	    RECT 0.6350 0.7300 0.8050 1.2450 ;
	    RECT 1.1450 0.7300 1.3150 2.0750 ;
	    RECT 2.9950 1.6550 3.1650 2.2450 ;
	    RECT 2.9950 1.2450 3.2550 1.6550 ;
	    RECT 0.5950 0.3200 0.8050 0.7300 ;
	    RECT 1.0950 0.3200 1.3150 0.7300 ;
   END
END efs8hd_and4b_2
MACRO efs8hd_and4bb_2
   CLASS CORE ;
   FOREIGN efs8hd_and4bb_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.6000 BY 3.4000 ;
   SITE unitehd ;
   PIN C
      PORT
         LAYER li1 ;
	    RECT 2.9050 0.5250 3.1750 1.6150 ;
      END
   END C
   PIN D
      PORT
         LAYER li1 ;
	    RECT 3.3500 0.5300 3.6550 1.7550 ;
      END
   END D
   PIN X
      PORT
         LAYER li1 ;
	    RECT 0.9900 1.9300 1.3200 2.1450 ;
	    RECT 1.0150 0.3200 1.2400 1.9300 ;
      END
   END X
   PIN BN
      PORT
         LAYER li1 ;
	    RECT 3.8250 0.7650 4.1750 1.6300 ;
      END
   END BN
   PIN AN
      PORT
         LAYER li1 ;
	    RECT 0.1450 1.1050 0.3300 2.0450 ;
      END
   END AN
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.4100 0.1050 1.7400 0.5800 ;
	    RECT 3.8350 0.1050 4.0050 0.5950 ;
	    RECT 0.5150 0.0850 4.0050 0.1050 ;
	    RECT 0.0000 -0.0850 4.6000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.6000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.6000 3.4850 ;
	    RECT 0.5150 3.2950 4.0850 3.3150 ;
	    RECT 0.5150 2.8200 0.8450 3.2950 ;
	    RECT 1.4900 2.8200 2.1600 3.2950 ;
	    RECT 2.7350 2.8200 3.0750 3.2950 ;
	    RECT 3.7550 2.8200 4.0850 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.6000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1750 2.5700 0.3450 3.0800 ;
	    RECT 2.3950 2.6050 2.5650 3.0800 ;
	    RECT 3.2450 2.6050 3.4150 3.0800 ;
	    RECT 4.2550 2.6050 4.5150 3.0800 ;
	    RECT 0.1750 2.3550 1.9250 2.5700 ;
	    RECT 0.5000 0.9350 0.6700 2.3550 ;
	    RECT 1.7550 1.6550 1.9250 2.3550 ;
	    RECT 2.2350 2.3950 3.4150 2.6050 ;
	    RECT 3.5850 2.3950 4.5150 2.6050 ;
	    RECT 0.1750 0.7650 0.6700 0.9350 ;
	    RECT 1.4150 1.0050 1.5850 1.6550 ;
	    RECT 1.7550 1.2450 2.0650 1.6550 ;
	    RECT 2.2350 1.0050 2.4050 2.3950 ;
	    RECT 3.5850 2.1800 3.7550 2.3950 ;
	    RECT 2.5750 1.9700 3.7550 2.1800 ;
	    RECT 2.5750 1.7500 2.7450 1.9700 ;
	    RECT 1.4150 0.7950 2.4050 1.0050 ;
	    RECT 0.1750 0.3200 0.3450 0.7650 ;
	    RECT 2.0100 0.3200 2.1800 0.7950 ;
	    RECT 4.3450 0.5950 4.5150 2.3950 ;
	    RECT 4.1750 0.3200 4.5150 0.5950 ;
   END
END efs8hd_and4bb_2
MACRO efs8hd_buf_12
   CLASS CORE ;
   FOREIGN efs8hd_buf_12 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 7.3600 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0950 0.1050 0.4250 0.7050 ;
	    RECT 0.9350 0.1050 1.2650 0.7050 ;
	    RECT 1.7750 0.1050 2.1050 0.7050 ;
	    RECT 2.6150 0.1050 2.9450 0.7050 ;
	    RECT 3.4550 0.1050 3.7850 0.7050 ;
	    RECT 4.2950 0.1050 4.6250 0.7050 ;
	    RECT 5.1350 0.1050 5.4650 0.7050 ;
	    RECT 5.9750 0.1050 6.3050 0.7050 ;
	    RECT 6.8150 0.1050 7.1450 1.1050 ;
	    RECT 0.0950 0.0850 7.1450 0.1050 ;
	    RECT 0.0000 -0.0850 7.3600 0.0850 ;
	    RECT 0.5700 -0.1050 0.7400 -0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 7.3600 0.3000 ;
      END
   END vgnd
   PIN X
      PORT
         LAYER li1 ;
	    RECT 2.2750 2.0200 2.4450 3.0800 ;
	    RECT 3.1150 2.0200 3.2850 3.0800 ;
	    RECT 3.9550 2.0200 4.1250 3.0800 ;
	    RECT 4.7950 2.0200 4.9650 3.0800 ;
	    RECT 5.6350 2.0200 5.8050 3.0800 ;
	    RECT 6.4750 2.0200 6.6450 3.0800 ;
	    RECT 2.2750 1.8050 6.6450 2.0200 ;
	    RECT 4.7100 1.1300 6.6450 1.8050 ;
	    RECT 2.2750 0.9200 6.6450 1.1300 ;
	    RECT 2.2750 0.3200 2.4450 0.9200 ;
	    RECT 3.1150 0.3200 3.2850 0.9200 ;
	    RECT 3.9550 0.3200 4.1250 0.9200 ;
	    RECT 4.7950 0.3200 4.9650 0.9200 ;
	    RECT 5.6350 0.3200 5.8050 0.9200 ;
	    RECT 6.4750 0.3200 6.6450 0.9200 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.1350 1.3450 1.6600 1.6150 ;
      END
   END A
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.5700 3.4850 0.7400 3.5050 ;
	    RECT 0.0000 3.3150 7.3600 3.4850 ;
	    RECT 0.1750 3.2950 7.1450 3.3150 ;
	    RECT 0.1750 2.2950 0.3450 3.2950 ;
	    RECT 1.0150 2.2950 1.1850 3.2950 ;
	    RECT 1.8550 2.2950 2.0250 3.2950 ;
	    RECT 2.6150 2.2950 2.9450 3.2950 ;
	    RECT 3.4550 2.2950 3.7850 3.2950 ;
	    RECT 4.2950 2.2950 4.6250 3.2950 ;
	    RECT 5.1350 2.2950 5.4650 3.2950 ;
	    RECT 5.9750 2.2950 6.3050 3.2950 ;
	    RECT 6.8150 1.8550 7.1450 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 7.3600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.5150 2.0200 0.8450 3.0800 ;
	    RECT 1.3550 2.0200 1.6850 3.0800 ;
	    RECT 0.5150 1.8050 2.0150 2.0200 ;
	    RECT 1.8400 1.5550 2.0150 1.8050 ;
	    RECT 1.8400 1.3450 4.4650 1.5550 ;
	    RECT 1.8400 1.1300 2.0150 1.3450 ;
	    RECT 0.5950 0.9200 2.0150 1.1300 ;
	    RECT 0.5950 0.3200 0.7650 0.9200 ;
	    RECT 1.4350 0.3250 1.6050 0.9200 ;
   END
END efs8hd_buf_12
MACRO efs8hd_buf_16
   CLASS CORE ;
   FOREIGN efs8hd_buf_16 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 10.1200 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3450 2.4850 1.6150 ;
      END
   END A
   PIN X
      PORT
         LAYER li1 ;
	    RECT 3.0350 2.0200 3.3650 3.0800 ;
	    RECT 3.8750 2.0200 4.2050 3.0800 ;
	    RECT 4.7150 2.0200 5.0450 3.0800 ;
	    RECT 5.5550 2.0200 5.8850 3.0800 ;
	    RECT 6.3950 2.0200 6.7250 3.0800 ;
	    RECT 7.2350 2.0200 7.5650 3.0800 ;
	    RECT 8.0750 2.0200 8.4050 3.0800 ;
	    RECT 8.9150 2.0200 9.2450 3.0800 ;
	    RECT 9.7600 2.0200 10.0350 2.9500 ;
	    RECT 3.0350 1.8050 10.0350 2.0200 ;
	    RECT 9.6550 1.1300 10.0350 1.8050 ;
	    RECT 3.0350 0.9200 10.0350 1.1300 ;
	    RECT 3.0350 0.3250 3.3650 0.9200 ;
	    RECT 3.8750 0.3250 4.2050 0.9200 ;
	    RECT 4.7150 0.3250 5.0450 0.9200 ;
	    RECT 5.5550 0.3250 5.8850 0.9200 ;
	    RECT 6.3950 0.3250 6.7250 0.9200 ;
	    RECT 7.2350 0.3250 7.5650 0.9200 ;
	    RECT 8.0750 0.3250 8.4050 0.9200 ;
	    RECT 8.9150 0.3250 9.2450 0.9200 ;
	    RECT 9.7600 0.4550 10.0350 0.9200 ;
	    RECT 3.0350 0.3200 3.2850 0.3250 ;
	    RECT 3.9550 0.3200 4.1250 0.3250 ;
	    RECT 4.7950 0.3200 4.9650 0.3250 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1750 0.1050 0.3450 1.1300 ;
	    RECT 1.0150 0.1050 1.1850 0.7050 ;
	    RECT 1.8550 0.1050 2.0250 0.7050 ;
	    RECT 2.6950 0.1050 2.8650 0.7050 ;
	    RECT 3.5350 0.1050 3.7050 0.7050 ;
	    RECT 4.3750 0.1050 4.5450 0.7050 ;
	    RECT 5.2150 0.1050 5.3850 0.7050 ;
	    RECT 6.0550 0.1050 6.2250 0.7050 ;
	    RECT 6.8950 0.1050 7.0650 0.7050 ;
	    RECT 7.7350 0.1050 7.9050 0.7050 ;
	    RECT 8.5750 0.1050 8.7450 0.7050 ;
	    RECT 9.4150 0.1050 9.5850 0.7050 ;
	    RECT 0.1750 0.0850 9.5850 0.1050 ;
	    RECT 0.0000 -0.0850 10.1200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 10.1200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 10.1200 3.4850 ;
	    RECT 0.1750 3.2950 9.5850 3.3150 ;
	    RECT 0.1750 1.8050 0.3450 3.2950 ;
	    RECT 1.0150 2.2950 1.1850 3.2950 ;
	    RECT 1.8550 2.2950 2.0250 3.2950 ;
	    RECT 2.6950 2.2950 2.8650 3.2950 ;
	    RECT 3.5350 2.2950 3.7050 3.2950 ;
	    RECT 4.3750 2.2950 4.5450 3.2950 ;
	    RECT 5.2150 2.2950 5.3850 3.2950 ;
	    RECT 6.0550 2.2950 6.2250 3.2950 ;
	    RECT 6.8950 2.2950 7.0650 3.2950 ;
	    RECT 7.7350 2.2950 7.9050 3.2950 ;
	    RECT 8.5750 2.2950 8.7450 3.2950 ;
	    RECT 9.4150 2.2950 9.5850 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 10.1200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.5150 2.0200 0.8450 3.0800 ;
	    RECT 1.3550 2.0200 1.6850 3.0800 ;
	    RECT 2.1950 2.0200 2.5250 3.0800 ;
	    RECT 0.5150 1.8050 2.8650 2.0200 ;
	    RECT 2.6900 1.5950 2.8650 1.8050 ;
	    RECT 2.6900 1.3450 9.4100 1.5950 ;
	    RECT 2.6900 1.1300 2.8650 1.3450 ;
	    RECT 0.5150 0.9200 2.8650 1.1300 ;
	    RECT 0.5150 0.3250 0.8450 0.9200 ;
	    RECT 1.3550 0.3250 1.6850 0.9200 ;
	    RECT 2.1950 0.3250 2.5250 0.9200 ;
   END
END efs8hd_buf_16
MACRO efs8hd_buf_2
   CLASS CORE ;
   FOREIGN efs8hd_buf_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 1.8400 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5600 0.1050 0.8900 0.5800 ;
	    RECT 1.4900 0.1050 1.7500 1.1550 ;
	    RECT 0.1450 0.0850 0.3150 0.1050 ;
	    RECT 0.5600 0.0850 1.7500 0.1050 ;
	    RECT 0.0000 -0.0850 1.8400 0.0850 ;
	    RECT 0.1450 -0.1050 0.3150 -0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 1.8400 0.3000 ;
      END
   END vgnd
   PIN X
      PORT
         LAYER li1 ;
	    RECT 1.0600 1.9500 1.3150 3.0800 ;
	    RECT 1.1450 1.0400 1.3150 1.9500 ;
	    RECT 1.0600 0.3200 1.3150 1.0400 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.1050 0.4400 1.6950 ;
      END
   END A
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.1450 3.4850 0.3150 3.5050 ;
	    RECT 0.0000 3.3150 1.8400 3.4850 ;
	    RECT 0.1450 3.2950 0.3150 3.3150 ;
	    RECT 0.5600 3.2950 1.7500 3.3150 ;
	    RECT 0.5600 2.3450 0.8900 3.2950 ;
	    RECT 1.4900 1.8550 1.7500 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 1.8400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1750 2.1300 0.3450 3.0800 ;
	    RECT 0.1750 1.9200 0.8900 2.1300 ;
	    RECT 0.7200 1.6550 0.8900 1.9200 ;
	    RECT 0.7200 1.2450 0.9750 1.6550 ;
	    RECT 0.7200 0.9350 0.8900 1.2450 ;
	    RECT 0.1750 0.7650 0.8900 0.9350 ;
	    RECT 0.1750 0.3200 0.3450 0.7650 ;
   END
END efs8hd_buf_2
MACRO efs8hd_buf_4
   CLASS CORE ;
   FOREIGN efs8hd_buf_4 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 2.7600 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5250 0.1050 0.7650 0.7050 ;
	    RECT 1.3550 0.1050 1.6850 0.7050 ;
	    RECT 2.1950 0.1050 2.5250 1.1050 ;
	    RECT 0.1500 0.0850 0.3200 0.1050 ;
	    RECT 0.5250 0.0850 2.5250 0.1050 ;
	    RECT 0.0000 -0.0850 2.7600 0.0850 ;
	    RECT 0.1500 -0.1050 0.3200 -0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 2.7600 0.3000 ;
      END
   END vgnd
   PIN X
      PORT
         LAYER li1 ;
	    RECT 1.0150 2.0200 1.1850 3.0800 ;
	    RECT 1.8550 2.0200 2.0250 3.0800 ;
	    RECT 1.0150 1.8050 2.0250 2.0200 ;
	    RECT 1.5250 1.1300 2.0250 1.8050 ;
	    RECT 1.0150 0.9200 2.0250 1.1300 ;
	    RECT 1.0150 0.3200 1.1850 0.9200 ;
	    RECT 1.8550 0.3200 2.0250 0.9200 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.3450 0.4700 1.6450 ;
      END
   END A
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.1500 3.4850 0.3200 3.5050 ;
	    RECT 0.0000 3.3150 2.7600 3.4850 ;
	    RECT 0.1500 3.2950 0.3200 3.3150 ;
	    RECT 0.5950 3.2950 2.5250 3.3150 ;
	    RECT 0.5950 2.2950 0.8350 3.2950 ;
	    RECT 1.3550 2.2950 1.6850 3.2950 ;
	    RECT 2.1950 1.8550 2.5250 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 2.7600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0950 2.0700 0.4250 3.0800 ;
	    RECT 0.0950 1.8550 0.8100 2.0700 ;
	    RECT 0.6400 1.5550 0.8100 1.8550 ;
	    RECT 0.6400 1.3450 1.1400 1.5550 ;
	    RECT 0.6400 1.1300 0.8100 1.3450 ;
	    RECT 0.1750 0.9200 0.8100 1.1300 ;
	    RECT 0.1750 0.3200 0.3450 0.9200 ;
   END
END efs8hd_buf_4
MACRO efs8hd_buf_6
   CLASS CORE ;
   FOREIGN efs8hd_buf_6 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.1400 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.4350 0.1050 0.6050 0.7050 ;
	    RECT 1.2750 0.1050 1.4450 0.7050 ;
	    RECT 2.0350 0.1050 2.3650 0.7050 ;
	    RECT 2.8750 0.1050 3.2050 0.7050 ;
	    RECT 3.7150 0.1050 4.0450 1.1050 ;
	    RECT 0.1500 0.0850 0.3200 0.1050 ;
	    RECT 0.4350 0.0850 4.0450 0.1050 ;
	    RECT 0.0000 -0.0850 4.1400 0.0850 ;
	    RECT 0.1500 -0.1050 0.3200 -0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.1400 0.3000 ;
      END
   END vgnd
   PIN X
      PORT
         LAYER li1 ;
	    RECT 1.6950 2.0200 1.8650 3.0800 ;
	    RECT 2.5350 2.0200 2.7050 3.0800 ;
	    RECT 3.3750 2.0200 3.5450 3.0800 ;
	    RECT 1.6950 1.8050 3.5450 2.0200 ;
	    RECT 2.2100 1.1300 3.5450 1.8050 ;
	    RECT 1.6950 0.9200 3.5450 1.1300 ;
	    RECT 1.6950 0.3200 1.8650 0.9200 ;
	    RECT 2.5350 0.3200 2.7050 0.9200 ;
	    RECT 3.3750 0.3200 3.5450 0.9200 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.1450 1.3450 1.1850 1.6450 ;
      END
   END A
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.1500 3.4850 0.3200 3.5050 ;
	    RECT 0.0000 3.3150 4.1400 3.4850 ;
	    RECT 0.1500 3.2950 0.3200 3.3150 ;
	    RECT 0.4350 3.2950 4.0450 3.3150 ;
	    RECT 0.4350 1.8550 0.6050 3.2950 ;
	    RECT 1.2750 2.2950 1.5150 3.2950 ;
	    RECT 2.0350 2.2950 2.3650 3.2950 ;
	    RECT 2.8750 2.2950 3.2050 3.2950 ;
	    RECT 3.7150 1.8550 4.0450 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.1400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.7750 2.0700 1.1050 3.0800 ;
	    RECT 0.7750 1.8550 1.5250 2.0700 ;
	    RECT 1.3550 1.5550 1.5250 1.8550 ;
	    RECT 1.3550 1.3450 1.8250 1.5550 ;
	    RECT 1.3550 1.1300 1.5250 1.3450 ;
	    RECT 0.7750 0.9200 1.5250 1.1300 ;
	    RECT 0.7750 0.3200 1.1050 0.9200 ;
   END
END efs8hd_buf_6
MACRO efs8hd_buf_8
   CLASS CORE ;
   FOREIGN efs8hd_buf_8 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.5200 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.7050 ;
	    RECT 1.3550 0.1050 1.6850 0.7050 ;
	    RECT 2.1950 0.1050 2.5250 0.7050 ;
	    RECT 3.0350 0.1050 3.3650 0.7050 ;
	    RECT 3.8750 0.1050 4.2050 0.7050 ;
	    RECT 4.7150 0.1050 5.0450 1.1050 ;
	    RECT 0.1500 0.0850 0.3200 0.1050 ;
	    RECT 0.5150 0.0850 5.0450 0.1050 ;
	    RECT 0.0000 -0.0850 5.5200 0.0850 ;
	    RECT 0.1500 -0.1050 0.3200 -0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.5200 0.3000 ;
      END
   END vgnd
   PIN X
      PORT
         LAYER li1 ;
	    RECT 1.8550 2.0200 2.0250 3.0800 ;
	    RECT 2.6950 2.0200 2.8650 3.0800 ;
	    RECT 3.5350 2.0200 3.7050 3.0800 ;
	    RECT 4.3750 2.0200 4.5450 3.0800 ;
	    RECT 1.8550 1.8050 4.5450 2.0200 ;
	    RECT 4.2850 1.1300 4.5450 1.8050 ;
	    RECT 1.8550 0.9200 4.5450 1.1300 ;
	    RECT 1.8550 0.3200 2.0250 0.9200 ;
	    RECT 2.6950 0.3200 2.8650 0.9200 ;
	    RECT 3.5350 0.3200 3.7050 0.9200 ;
	    RECT 4.3750 0.3200 4.5450 0.9200 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.1400 1.3450 1.2400 1.6150 ;
      END
   END A
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.1500 3.4850 0.3200 3.5050 ;
	    RECT 0.0000 3.3150 5.5200 3.4850 ;
	    RECT 0.1500 3.2950 0.3200 3.3150 ;
	    RECT 0.5950 3.2950 5.0450 3.3150 ;
	    RECT 0.5950 2.2950 0.7650 3.2950 ;
	    RECT 1.4350 2.2950 1.6050 3.2950 ;
	    RECT 2.1950 2.2950 2.5250 3.2950 ;
	    RECT 3.0350 2.2950 3.3650 3.2950 ;
	    RECT 3.8750 2.2950 4.2050 3.2950 ;
	    RECT 4.7150 1.8550 5.0450 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.5200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0950 2.0200 0.4250 3.0800 ;
	    RECT 0.9350 2.0200 1.2650 3.0800 ;
	    RECT 0.0950 1.8050 1.5950 2.0200 ;
	    RECT 1.4200 1.5550 1.5950 1.8050 ;
	    RECT 1.4200 1.3450 4.0450 1.5550 ;
	    RECT 1.4200 1.1300 1.5950 1.3450 ;
	    RECT 0.1750 0.9200 1.5950 1.1300 ;
	    RECT 0.1750 0.3200 0.3450 0.9200 ;
	    RECT 1.0150 0.3250 1.1850 0.9200 ;
   END
END efs8hd_buf_8
MACRO efs8hd_bufbuf_16
   CLASS CORE ;
   FOREIGN efs8hd_bufbuf_16 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 11.9600 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.1100 1.3450 0.4400 1.6150 ;
      END
   END A
   PIN X
      PORT
         LAYER li1 ;
	    RECT 5.2350 2.0200 5.5650 3.0800 ;
	    RECT 6.0750 2.0200 6.4050 3.0800 ;
	    RECT 6.9150 2.0200 7.2450 3.0800 ;
	    RECT 7.7550 2.0200 8.0850 3.0800 ;
	    RECT 8.5950 2.0200 8.9250 3.0800 ;
	    RECT 9.4350 2.0200 9.7650 3.0800 ;
	    RECT 10.2750 2.0200 10.6050 3.0800 ;
	    RECT 11.1150 2.0200 11.4450 3.0800 ;
	    RECT 5.2350 1.8050 11.8750 2.0200 ;
	    RECT 11.6200 1.1300 11.8750 1.8050 ;
	    RECT 5.2350 0.9200 11.8750 1.1300 ;
	    RECT 5.2350 0.3250 5.5650 0.9200 ;
	    RECT 6.0750 0.3250 6.4050 0.9200 ;
	    RECT 6.9150 0.3250 7.2450 0.9200 ;
	    RECT 7.7550 0.3250 8.0850 0.9200 ;
	    RECT 8.5950 0.3250 8.9250 0.9200 ;
	    RECT 9.4350 0.3250 9.7650 0.9200 ;
	    RECT 10.2750 0.3250 10.6050 0.9200 ;
	    RECT 11.1150 0.3250 11.4450 0.9200 ;
	    RECT 5.2350 0.3200 5.4850 0.3250 ;
	    RECT 6.1550 0.3200 6.3250 0.3250 ;
	    RECT 6.9950 0.3200 7.1650 0.3250 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1750 0.1050 0.3450 1.1300 ;
	    RECT 1.5350 0.1050 1.7050 0.7050 ;
	    RECT 2.3750 0.1050 2.5450 0.7050 ;
	    RECT 3.2150 0.1050 3.3850 0.7050 ;
	    RECT 4.0550 0.1050 4.2250 0.7050 ;
	    RECT 4.8950 0.1050 5.0650 0.7050 ;
	    RECT 5.7350 0.1050 5.9050 0.7050 ;
	    RECT 6.5750 0.1050 6.7450 0.7050 ;
	    RECT 7.4150 0.1050 7.5850 0.7050 ;
	    RECT 8.2550 0.1050 8.4250 0.7050 ;
	    RECT 9.0950 0.1050 9.2650 0.7050 ;
	    RECT 9.9350 0.1050 10.1050 0.7050 ;
	    RECT 10.7750 0.1050 10.9450 0.7050 ;
	    RECT 11.6150 0.1050 11.7850 0.7050 ;
	    RECT 0.1750 0.0850 11.7850 0.1050 ;
	    RECT 0.0000 -0.0850 11.9600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 11.9600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 11.9600 3.4850 ;
	    RECT 0.1750 3.2950 11.7850 3.3150 ;
	    RECT 0.1750 1.8050 0.3450 3.2950 ;
	    RECT 1.5350 2.2300 1.7050 3.2950 ;
	    RECT 2.3750 2.2300 2.5450 3.2950 ;
	    RECT 3.2150 2.2950 3.3850 3.2950 ;
	    RECT 4.0550 2.2950 4.2250 3.2950 ;
	    RECT 4.8950 2.2950 5.0650 3.2950 ;
	    RECT 5.7350 2.2950 5.9050 3.2950 ;
	    RECT 6.5750 2.2950 6.7450 3.2950 ;
	    RECT 7.4150 2.2950 7.5850 3.2950 ;
	    RECT 8.2550 2.2950 8.4250 3.2950 ;
	    RECT 9.0950 2.2950 9.2650 3.2950 ;
	    RECT 9.9350 2.2950 10.1050 3.2950 ;
	    RECT 10.7750 2.2950 10.9450 3.2950 ;
	    RECT 11.6150 2.2950 11.7850 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 11.9600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.5150 1.8050 0.8450 3.0800 ;
	    RECT 1.0350 2.0200 1.3650 3.0800 ;
	    RECT 1.8750 2.0200 2.2050 3.0800 ;
	    RECT 2.7150 2.0200 3.0450 3.0800 ;
	    RECT 3.5550 2.0200 3.8850 3.0800 ;
	    RECT 4.3950 2.0200 4.7250 3.0800 ;
	    RECT 1.0350 1.8050 2.5450 2.0200 ;
	    RECT 2.7150 1.8050 5.0650 2.0200 ;
	    RECT 0.6100 1.5950 0.8450 1.8050 ;
	    RECT 2.3750 1.5950 2.5450 1.8050 ;
	    RECT 4.8900 1.5950 5.0650 1.8050 ;
	    RECT 0.6100 1.3450 2.2050 1.5950 ;
	    RECT 2.3750 1.3450 4.6850 1.5950 ;
	    RECT 4.8900 1.3450 11.4500 1.5950 ;
	    RECT 0.6100 1.1300 0.8450 1.3450 ;
	    RECT 2.3750 1.1300 2.5450 1.3450 ;
	    RECT 4.8900 1.1300 5.0650 1.3450 ;
	    RECT 0.5150 0.3250 0.8450 1.1300 ;
	    RECT 1.0350 0.9200 2.5450 1.1300 ;
	    RECT 2.7150 0.9200 5.0650 1.1300 ;
	    RECT 1.0350 0.3250 1.3650 0.9200 ;
	    RECT 1.8750 0.3250 2.2050 0.9200 ;
	    RECT 2.7150 0.3250 3.0450 0.9200 ;
	    RECT 3.5550 0.3250 3.8850 0.9200 ;
	    RECT 4.3950 0.3250 4.7250 0.9200 ;
   END
END efs8hd_bufbuf_16
MACRO efs8hd_bufbuf_8
   CLASS CORE ;
   FOREIGN efs8hd_bufbuf_8 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 6.9000 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.1100 1.3450 0.4400 1.6150 ;
      END
   END A
   PIN X
      PORT
         LAYER li1 ;
	    RECT 3.2300 2.0200 3.5600 3.0800 ;
	    RECT 4.0700 2.0200 4.4000 3.0800 ;
	    RECT 4.9100 2.0200 5.2400 3.0800 ;
	    RECT 5.7500 2.0200 6.0800 3.0800 ;
	    RECT 3.2300 1.8050 6.8150 2.0200 ;
	    RECT 6.4350 1.1300 6.8150 1.8050 ;
	    RECT 3.2300 0.9200 6.8150 1.1300 ;
	    RECT 3.2300 0.3250 3.5600 0.9200 ;
	    RECT 4.0700 0.3250 4.4000 0.9200 ;
	    RECT 4.9100 0.3250 5.2400 0.9200 ;
	    RECT 5.7500 0.3250 6.0800 0.9200 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5950 0.1050 0.7650 0.7050 ;
	    RECT 2.0500 0.1050 2.2200 0.7050 ;
	    RECT 2.8900 0.1050 3.0600 0.7050 ;
	    RECT 3.7300 0.1050 3.9000 0.7050 ;
	    RECT 4.5700 0.1050 4.7400 0.7050 ;
	    RECT 5.4100 0.1050 5.5800 0.7050 ;
	    RECT 6.2500 0.1050 6.4200 0.7050 ;
	    RECT 0.5950 0.0850 6.4200 0.1050 ;
	    RECT 0.0000 -0.0850 6.9000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 6.9000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 6.9000 3.4850 ;
	    RECT 0.5950 3.2950 6.4200 3.3150 ;
	    RECT 0.5950 2.2300 0.7650 3.2950 ;
	    RECT 2.0500 2.2300 2.2200 3.2950 ;
	    RECT 2.8900 2.2300 3.0600 3.2950 ;
	    RECT 3.7300 2.2950 3.9000 3.2950 ;
	    RECT 4.5700 2.2950 4.7400 3.2950 ;
	    RECT 5.4100 2.2950 5.5800 3.2950 ;
	    RECT 6.2500 2.2950 6.4200 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 6.9000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0950 2.0200 0.4250 2.7000 ;
	    RECT 0.0950 1.8050 0.7800 2.0200 ;
	    RECT 1.0000 1.9300 1.3800 3.0800 ;
	    RECT 0.6100 1.6550 0.7800 1.8050 ;
	    RECT 0.6100 1.2450 1.0400 1.6550 ;
	    RECT 1.2100 1.5950 1.3800 1.9300 ;
	    RECT 1.5500 2.0200 1.8800 3.0800 ;
	    RECT 2.3900 2.0200 2.7200 3.0800 ;
	    RECT 1.5500 1.8050 3.0600 2.0200 ;
	    RECT 2.8900 1.5950 3.0600 1.8050 ;
	    RECT 1.2100 1.3450 2.7200 1.5950 ;
	    RECT 2.8900 1.3450 5.3600 1.5950 ;
	    RECT 0.6100 1.1300 0.7800 1.2450 ;
	    RECT 0.0950 0.9200 0.7800 1.1300 ;
	    RECT 1.2100 1.0300 1.3800 1.3450 ;
	    RECT 2.8900 1.1300 3.0600 1.3450 ;
	    RECT 0.0950 0.3250 0.4250 0.9200 ;
	    RECT 1.0000 0.3250 1.3800 1.0300 ;
	    RECT 1.5500 0.9200 3.0600 1.1300 ;
	    RECT 1.5500 0.3250 1.8800 0.9200 ;
	    RECT 2.3900 0.3250 2.7200 0.9200 ;
   END
END efs8hd_bufbuf_8
MACRO efs8hd_bufinv_16
   CLASS CORE ;
   FOREIGN efs8hd_bufinv_16 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 11.0400 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.3450 1.2650 1.6150 ;
      END
   END A
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 4.2950 2.0200 4.6250 3.0800 ;
	    RECT 5.1350 2.0200 5.4650 3.0800 ;
	    RECT 5.9750 2.0200 6.3050 3.0800 ;
	    RECT 6.8150 2.0200 7.1450 3.0800 ;
	    RECT 7.6550 2.0200 7.9850 3.0800 ;
	    RECT 8.4950 2.0200 8.8250 3.0800 ;
	    RECT 9.3350 2.0200 9.6650 3.0800 ;
	    RECT 10.1750 2.0200 10.5050 3.0800 ;
	    RECT 4.2950 1.8050 10.9550 2.0200 ;
	    RECT 10.6800 1.1300 10.9550 1.8050 ;
	    RECT 4.2950 0.9200 10.9550 1.1300 ;
	    RECT 4.2950 0.3250 4.6250 0.9200 ;
	    RECT 5.1350 0.3250 5.4650 0.9200 ;
	    RECT 5.9750 0.3250 6.3050 0.9200 ;
	    RECT 6.8150 0.3250 7.1450 0.9200 ;
	    RECT 7.6550 0.3250 7.9850 0.9200 ;
	    RECT 8.4950 0.3250 8.8250 0.9200 ;
	    RECT 9.3350 0.3250 9.6650 0.9200 ;
	    RECT 10.1750 0.3250 10.5050 0.9200 ;
	    RECT 4.2950 0.3200 4.5450 0.3250 ;
	    RECT 5.2150 0.3200 5.3850 0.3250 ;
	    RECT 6.0550 0.3200 6.2250 0.3250 ;
      END
   END Y
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5950 0.1050 0.7650 0.7050 ;
	    RECT 1.4350 0.1050 1.6050 0.7050 ;
	    RECT 2.2750 0.1050 2.4450 0.7050 ;
	    RECT 3.1150 0.1050 3.2850 0.7050 ;
	    RECT 3.9550 0.1050 4.1250 0.7050 ;
	    RECT 4.7950 0.1050 4.9650 0.7050 ;
	    RECT 5.6350 0.1050 5.8050 0.7050 ;
	    RECT 6.4750 0.1050 6.6450 0.7050 ;
	    RECT 7.3150 0.1050 7.4850 0.7050 ;
	    RECT 8.1550 0.1050 8.3250 0.7050 ;
	    RECT 8.9950 0.1050 9.1650 0.7050 ;
	    RECT 9.8350 0.1050 10.0050 0.7050 ;
	    RECT 10.6750 0.1050 10.8450 0.7050 ;
	    RECT 0.5950 0.0850 10.8450 0.1050 ;
	    RECT 0.0000 -0.0850 11.0400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 11.0400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 11.0400 3.4850 ;
	    RECT 0.5950 3.2950 10.8450 3.3150 ;
	    RECT 0.5950 2.2300 0.7650 3.2950 ;
	    RECT 1.4350 2.2300 1.6050 3.2950 ;
	    RECT 2.2750 2.2950 2.4450 3.2950 ;
	    RECT 3.1150 2.2950 3.2850 3.2950 ;
	    RECT 3.9550 2.2950 4.1250 3.2950 ;
	    RECT 4.7950 2.2950 4.9650 3.2950 ;
	    RECT 5.6350 2.2950 5.8050 3.2950 ;
	    RECT 6.4750 2.2950 6.6450 3.2950 ;
	    RECT 7.3150 2.2950 7.4850 3.2950 ;
	    RECT 8.1550 2.2950 8.3250 3.2950 ;
	    RECT 8.9950 2.2950 9.1650 3.2950 ;
	    RECT 9.8350 2.2950 10.0050 3.2950 ;
	    RECT 10.6750 2.2950 10.8450 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 11.0400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0950 2.0200 0.4250 3.0800 ;
	    RECT 0.9350 2.0200 1.2650 3.0800 ;
	    RECT 1.7750 2.0200 2.1050 3.0800 ;
	    RECT 2.6150 2.0200 2.9450 3.0800 ;
	    RECT 3.4550 2.0200 3.7850 3.0800 ;
	    RECT 0.0950 1.8050 1.6050 2.0200 ;
	    RECT 1.7750 1.8050 4.1250 2.0200 ;
	    RECT 1.4350 1.5950 1.6050 1.8050 ;
	    RECT 3.9500 1.5950 4.1250 1.8050 ;
	    RECT 1.4350 1.3450 3.7450 1.5950 ;
	    RECT 3.9500 1.3450 10.5100 1.5950 ;
	    RECT 1.4350 1.1300 1.6050 1.3450 ;
	    RECT 3.9500 1.1300 4.1250 1.3450 ;
	    RECT 0.0950 0.9200 1.6050 1.1300 ;
	    RECT 1.7750 0.9200 4.1250 1.1300 ;
	    RECT 0.0950 0.3250 0.4250 0.9200 ;
	    RECT 0.9350 0.3250 1.2650 0.9200 ;
	    RECT 1.7750 0.3250 2.1050 0.9200 ;
	    RECT 2.6150 0.3250 2.9450 0.9200 ;
	    RECT 3.4550 0.3250 3.7850 0.9200 ;
   END
END efs8hd_bufinv_16
MACRO efs8hd_bufinv_8
   CLASS CORE ;
   FOREIGN efs8hd_bufinv_8 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 6.4400 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3450 0.5050 1.6150 ;
      END
   END A
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 2.7150 2.0200 3.0450 3.0800 ;
	    RECT 3.5550 2.0200 3.8850 3.0800 ;
	    RECT 4.3950 2.0200 4.7250 3.0800 ;
	    RECT 5.2350 2.0200 5.5650 3.0800 ;
	    RECT 2.7150 1.8050 6.3550 2.0200 ;
	    RECT 5.9700 1.1300 6.3550 1.8050 ;
	    RECT 2.7150 0.9200 6.3550 1.1300 ;
	    RECT 2.7150 0.3250 3.0450 0.9200 ;
	    RECT 3.5550 0.3250 3.8850 0.9200 ;
	    RECT 4.3950 0.3250 4.7250 0.9200 ;
	    RECT 5.2350 0.3250 5.5650 0.9200 ;
      END
   END Y
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1750 0.1050 0.3450 1.1300 ;
	    RECT 1.5350 0.1050 1.7050 0.7050 ;
	    RECT 2.3750 0.1050 2.5450 0.7050 ;
	    RECT 3.2150 0.1050 3.3850 0.7050 ;
	    RECT 4.0550 0.1050 4.2250 0.7050 ;
	    RECT 4.8950 0.1050 5.0650 0.7050 ;
	    RECT 5.7350 0.1050 5.9050 0.7050 ;
	    RECT 0.1750 0.0850 5.9050 0.1050 ;
	    RECT 0.0000 -0.0850 6.4400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 6.4400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 6.4400 3.4850 ;
	    RECT 0.1750 3.2950 5.9050 3.3150 ;
	    RECT 0.1750 1.8050 0.3450 3.2950 ;
	    RECT 1.5350 2.2300 1.7050 3.2950 ;
	    RECT 2.3750 2.2300 2.5450 3.2950 ;
	    RECT 3.2150 2.2950 3.3850 3.2950 ;
	    RECT 4.0550 2.2950 4.2250 3.2950 ;
	    RECT 4.8950 2.2950 5.0650 3.2950 ;
	    RECT 5.7350 2.2950 5.9050 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 6.4400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.5150 1.9300 0.8450 3.0800 ;
	    RECT 0.6750 1.5950 0.8450 1.9300 ;
	    RECT 1.0350 2.0200 1.3650 3.0800 ;
	    RECT 1.8750 2.0200 2.2050 3.0800 ;
	    RECT 1.0350 1.8050 2.5450 2.0200 ;
	    RECT 2.3750 1.5950 2.5450 1.8050 ;
	    RECT 0.6750 1.3450 2.2050 1.5950 ;
	    RECT 2.3750 1.3450 5.7600 1.5950 ;
	    RECT 0.6750 1.1300 0.8450 1.3450 ;
	    RECT 2.3750 1.1300 2.5450 1.3450 ;
	    RECT 0.5150 0.3250 0.8450 1.1300 ;
	    RECT 1.0350 0.9200 2.5450 1.1300 ;
	    RECT 1.0350 0.3250 1.3650 0.9200 ;
	    RECT 1.8750 0.3250 2.2050 0.9200 ;
   END
END efs8hd_bufinv_8
MACRO efs8hd_clkbuf_16
   CLASS CORE ;
   FOREIGN efs8hd_clkbuf_16 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 9.2000 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.7650 0.4000 1.6550 ;
      END
   END A
   PIN X
      PORT
         LAYER li1 ;
	    RECT 2.2800 2.1700 2.5400 3.0750 ;
	    RECT 3.1400 2.1700 3.4000 3.0750 ;
	    RECT 4.0000 2.1700 4.2600 3.0750 ;
	    RECT 4.8600 2.1700 5.1200 3.0750 ;
	    RECT 5.7050 2.1700 5.9650 3.0750 ;
	    RECT 6.5650 2.1700 6.8250 3.0750 ;
	    RECT 7.4250 2.1700 7.6850 3.0750 ;
	    RECT 2.2800 2.1500 7.6850 2.1700 ;
	    RECT 8.2950 2.1500 8.5850 3.0750 ;
	    RECT 2.2800 1.8700 9.0250 2.1500 ;
	    RECT 7.8600 1.1300 9.0250 1.8700 ;
	    RECT 2.2800 0.9200 9.0250 1.1300 ;
	    RECT 2.2800 0.3500 2.5400 0.9200 ;
	    RECT 3.1400 0.3500 3.4000 0.9200 ;
	    RECT 4.0000 0.3500 4.2600 0.9200 ;
	    RECT 4.8450 0.3500 5.1200 0.9200 ;
	    RECT 5.7050 0.3500 5.9650 0.9200 ;
	    RECT 6.5650 0.3500 6.8250 0.9200 ;
	    RECT 7.4250 0.3500 7.6850 0.9200 ;
	    RECT 8.2950 0.3500 8.5550 0.9200 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.1050 0.4250 0.5950 ;
	    RECT 0.9900 0.1050 1.2500 0.7650 ;
	    RECT 1.8500 0.1050 2.1100 0.8050 ;
	    RECT 2.7100 0.1050 2.9700 0.7050 ;
	    RECT 3.5700 0.1050 3.8300 0.7050 ;
	    RECT 4.4300 0.1050 4.6750 0.7050 ;
	    RECT 5.2900 0.1050 5.5350 0.7050 ;
	    RECT 6.1450 0.1050 6.3950 0.7050 ;
	    RECT 7.0050 0.1050 7.2550 0.7050 ;
	    RECT 7.8650 0.1050 8.1250 0.7050 ;
	    RECT 8.7250 0.1050 9.0250 0.7050 ;
	    RECT 0.0850 0.0850 9.0250 0.1050 ;
	    RECT 0.0000 -0.0850 9.2000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 9.2000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 9.2000 3.4850 ;
	    RECT 0.0950 3.2950 9.0250 3.3150 ;
	    RECT 0.0950 2.2800 0.3900 3.2950 ;
	    RECT 0.9900 2.2800 1.2500 3.2950 ;
	    RECT 1.8500 3.2900 8.1250 3.2950 ;
	    RECT 1.8500 2.2950 2.1100 3.2900 ;
	    RECT 2.7100 2.3800 2.9700 3.2900 ;
	    RECT 3.5700 2.3800 3.8300 3.2900 ;
	    RECT 4.4300 2.3800 4.6900 3.2900 ;
	    RECT 5.2900 2.3800 5.5350 3.2900 ;
	    RECT 6.1500 2.3800 6.3950 3.2900 ;
	    RECT 7.0100 2.3800 7.2550 3.2900 ;
	    RECT 7.8700 2.3800 8.1250 3.2900 ;
	    RECT 8.7550 2.3650 9.0250 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 9.2000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.5950 1.6550 0.8150 3.0800 ;
	    RECT 1.4300 1.6550 1.6800 3.0750 ;
	    RECT 0.5950 1.3450 7.6900 1.6550 ;
	    RECT 0.5950 0.3300 0.8200 1.3450 ;
	    RECT 1.4300 0.3300 1.6800 1.3450 ;
   END
END efs8hd_clkbuf_16
MACRO efs8hd_clkbuf_2
   CLASS CORE ;
   FOREIGN efs8hd_clkbuf_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 1.8400 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.4450 0.7650 0.7850 1.6550 ;
      END
   END A
   PIN X
      PORT
         LAYER li1 ;
	    RECT 1.0600 2.5400 1.2450 3.0450 ;
	    RECT 1.0600 2.3200 1.7250 2.5400 ;
	    RECT 1.3850 1.0300 1.7250 2.3200 ;
	    RECT 1.0400 0.8200 1.7250 1.0300 ;
	    RECT 1.0400 0.3200 1.2450 0.8200 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5250 0.1050 0.8550 0.5950 ;
	    RECT 1.4150 0.1050 1.7500 0.6050 ;
	    RECT 0.5250 0.0850 1.7500 0.1050 ;
	    RECT 0.0000 -0.0850 1.8400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 1.8400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 1.8400 3.4850 ;
	    RECT 0.5250 3.2950 1.7500 3.3150 ;
	    RECT 0.5250 2.3200 0.8550 3.2950 ;
	    RECT 1.4150 2.7650 1.7500 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 1.8400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.0800 0.3550 3.0450 ;
	    RECT 0.0850 1.8700 1.2150 2.0800 ;
	    RECT 0.0850 0.6250 0.2550 1.8700 ;
	    RECT 0.9650 1.2450 1.2150 1.8700 ;
	    RECT 0.0850 0.2950 0.3450 0.6250 ;
   END
END efs8hd_clkbuf_2
MACRO efs8hd_clkbuf_4
   CLASS CORE ;
   FOREIGN efs8hd_clkbuf_4 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 2.7600 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.4250 0.7650 0.7750 1.6550 ;
      END
   END A
   PIN X
      PORT
         LAYER li1 ;
	    RECT 1.0450 2.5050 1.3050 3.0800 ;
	    RECT 1.9050 2.5050 2.1650 3.0800 ;
	    RECT 1.0450 2.2950 2.1650 2.5050 ;
	    RECT 1.9050 1.9800 2.1650 2.2950 ;
	    RECT 1.9050 1.7700 2.6600 1.9800 ;
	    RECT 2.2550 1.1300 2.6600 1.7700 ;
	    RECT 1.0100 0.9200 2.6600 1.1300 ;
	    RECT 1.0100 0.4300 1.3050 0.9200 ;
	    RECT 1.9050 0.4300 2.1650 0.9200 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5950 0.1050 0.8300 0.5950 ;
	    RECT 1.4750 0.1050 1.7300 0.7050 ;
	    RECT 2.3350 0.1050 2.6150 0.7050 ;
	    RECT 0.5950 0.0850 2.6150 0.1050 ;
	    RECT 0.0000 -0.0850 2.7600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 2.7600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 2.7600 3.4850 ;
	    RECT 0.5650 3.2950 2.6200 3.3150 ;
	    RECT 0.5650 2.2950 0.8750 3.2950 ;
	    RECT 1.4750 2.7200 1.7300 3.2950 ;
	    RECT 2.3350 2.2050 2.6200 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 2.7600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.0800 0.3950 3.0800 ;
	    RECT 0.0850 1.8700 1.1150 2.0800 ;
	    RECT 0.0850 0.5950 0.2550 1.8700 ;
	    RECT 0.9450 1.5550 1.1150 1.8700 ;
	    RECT 0.9450 1.3450 2.0850 1.5550 ;
	    RECT 0.0850 0.3200 0.4250 0.5950 ;
   END
END efs8hd_clkbuf_4
MACRO efs8hd_clkbuf_8
   CLASS CORE ;
   FOREIGN efs8hd_clkbuf_8 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.0600 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.7650 0.4000 1.6550 ;
      END
   END A
   PIN X
      PORT
         LAYER li1 ;
	    RECT 1.4200 2.1700 1.6800 3.0750 ;
	    RECT 2.2800 2.1700 2.5400 3.0750 ;
	    RECT 3.1400 2.1700 3.4000 3.0750 ;
	    RECT 4.0000 2.1700 4.2600 3.0750 ;
	    RECT 1.4200 1.8700 4.7300 2.1700 ;
	    RECT 3.7600 1.1300 4.7300 1.8700 ;
	    RECT 1.4200 0.9200 4.7300 1.1300 ;
	    RECT 1.4200 0.3500 1.6800 0.9200 ;
	    RECT 2.2800 0.3500 2.5400 0.9200 ;
	    RECT 3.1400 0.3500 3.4000 0.9200 ;
	    RECT 4.0000 0.3500 4.2600 0.9200 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1450 0.1050 0.3900 0.5950 ;
	    RECT 0.9900 0.1050 1.2500 0.7650 ;
	    RECT 1.8500 0.1050 2.1100 0.7050 ;
	    RECT 2.7100 0.1050 2.9700 0.7050 ;
	    RECT 3.5700 0.1050 3.8300 0.7050 ;
	    RECT 4.4300 0.1050 4.7300 0.7050 ;
	    RECT 0.1450 0.0850 4.7300 0.1050 ;
	    RECT 0.0000 -0.0850 5.0600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.0600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.0600 3.4850 ;
	    RECT 0.0950 3.2950 4.7250 3.3150 ;
	    RECT 0.0950 1.9050 0.3900 3.2950 ;
	    RECT 0.9900 1.9050 1.2500 3.2950 ;
	    RECT 1.8500 2.3800 2.1100 3.2950 ;
	    RECT 2.7100 2.3800 2.9700 3.2950 ;
	    RECT 3.5700 2.3800 3.8300 3.2950 ;
	    RECT 4.4300 2.3800 4.7250 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.0600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.5700 1.6550 0.8200 3.0750 ;
	    RECT 0.5700 1.3450 3.5900 1.6550 ;
	    RECT 0.5700 0.3300 0.8200 1.3450 ;
   END
END efs8hd_clkbuf_8
MACRO efs8hd_clkdlybuf4s15_1
   CLASS CORE ;
   FOREIGN efs8hd_clkdlybuf4s15_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.6800 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 3.2100 2.2000 3.5950 3.0800 ;
	    RECT 3.3650 0.6800 3.5950 2.2000 ;
	    RECT 3.2100 0.3550 3.5950 0.6800 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3200 0.5600 1.6550 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5950 0.1050 0.9100 0.6800 ;
	    RECT 2.7100 0.1050 3.0400 0.6800 ;
	    RECT 0.5950 0.0850 3.0400 0.1050 ;
	    RECT 0.0000 -0.0850 3.6800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.6800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.6800 3.4850 ;
	    RECT 0.5950 3.2950 3.0400 3.3150 ;
	    RECT 0.5950 2.2950 0.9250 3.2950 ;
	    RECT 2.6400 2.2000 3.0400 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.6800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.0800 0.4250 3.0800 ;
	    RECT 1.3850 2.2950 1.7600 3.0800 ;
	    RECT 0.0850 1.8700 1.2150 2.0800 ;
	    RECT 0.7300 1.1050 1.2150 1.8700 ;
	    RECT 0.0850 0.8950 1.2150 1.1050 ;
	    RECT 1.5900 1.5650 1.7600 2.2950 ;
	    RECT 1.9300 1.9900 2.4100 3.0800 ;
	    RECT 1.9300 1.7750 3.1950 1.9900 ;
	    RECT 1.5900 1.3200 2.6850 1.5650 ;
	    RECT 1.5900 1.0300 1.7600 1.3200 ;
	    RECT 2.8550 1.1050 3.1950 1.7750 ;
	    RECT 0.0850 0.3200 0.4250 0.8950 ;
	    RECT 1.3850 0.3200 1.7600 1.0300 ;
	    RECT 1.9300 0.8950 3.1950 1.1050 ;
	    RECT 1.9300 0.3200 2.2600 0.8950 ;
   END
END efs8hd_clkdlybuf4s15_1
MACRO efs8hd_clkdlybuf4s15_2
   CLASS CORE ;
   FOREIGN efs8hd_clkdlybuf4s15_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.1400 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 3.0700 1.8550 3.5500 3.0800 ;
	    RECT 3.3550 0.8000 3.5500 1.8550 ;
	    RECT 3.0500 0.3200 3.5500 0.8000 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3250 0.5550 2.0300 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5850 0.1050 0.9150 0.6900 ;
	    RECT 2.5500 0.1050 2.8800 0.7050 ;
	    RECT 3.7200 0.1050 4.0550 0.8050 ;
	    RECT 0.5850 0.0850 4.0550 0.1050 ;
	    RECT 0.0000 -0.0850 4.1400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.1400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.1400 3.4850 ;
	    RECT 0.6000 3.2950 4.0550 3.3150 ;
	    RECT 0.6000 2.6700 0.9300 3.2950 ;
	    RECT 2.5500 2.6700 2.8800 3.2950 ;
	    RECT 3.7200 1.8550 4.0550 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.1400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.4550 0.4300 3.0800 ;
	    RECT 0.0850 2.2450 1.0600 2.4550 ;
	    RECT 0.8900 1.5550 1.0600 2.2450 ;
	    RECT 1.2300 2.2300 1.6600 3.0800 ;
	    RECT 1.8300 2.4550 2.1000 3.0800 ;
	    RECT 1.8300 2.2400 2.9000 2.4550 ;
	    RECT 1.4900 1.8550 1.6600 2.2300 ;
	    RECT 0.8900 1.3450 1.3200 1.5550 ;
	    RECT 1.4900 1.3450 2.4150 1.8550 ;
	    RECT 2.7300 1.5550 2.9000 2.2400 ;
	    RECT 2.7300 1.3450 3.1850 1.5550 ;
	    RECT 0.8900 1.1150 1.0600 1.3450 ;
	    RECT 1.4900 1.1300 1.6600 1.3450 ;
	    RECT 2.7300 1.1300 2.9000 1.3450 ;
	    RECT 0.0850 0.9000 1.0600 1.1150 ;
	    RECT 0.0850 0.3200 0.4150 0.9000 ;
	    RECT 1.2800 0.3200 1.6600 1.1300 ;
	    RECT 1.8300 0.9200 2.9000 1.1300 ;
	    RECT 1.8300 0.3200 2.1000 0.9200 ;
   END
END efs8hd_clkdlybuf4s15_2
MACRO efs8hd_clkdlybuf4s18_1
   CLASS CORE ;
   FOREIGN efs8hd_clkdlybuf4s18_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.6800 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 3.2200 2.2000 3.5900 3.0800 ;
	    RECT 3.3650 0.6800 3.5900 2.2000 ;
	    RECT 3.2100 0.3200 3.5900 0.6800 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.1000 1.3200 0.5500 1.6550 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5950 0.1050 0.9100 0.6800 ;
	    RECT 2.7100 0.1050 3.0400 0.6800 ;
	    RECT 0.5950 0.0850 3.0400 0.1050 ;
	    RECT 0.0000 -0.0850 3.6800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.6800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.6800 3.4850 ;
	    RECT 0.5950 3.2950 3.0400 3.3150 ;
	    RECT 0.5950 2.2950 0.9250 3.2950 ;
	    RECT 2.7100 2.2000 3.0400 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.6800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0950 2.0800 0.4250 3.0800 ;
	    RECT 1.3850 2.2950 1.7600 3.0800 ;
	    RECT 0.0950 1.8700 1.2150 2.0800 ;
	    RECT 0.7200 1.1050 1.2150 1.8700 ;
	    RECT 0.0950 0.8950 1.2150 1.1050 ;
	    RECT 1.5900 1.5650 1.7600 2.2950 ;
	    RECT 1.9300 1.9900 2.2600 3.0800 ;
	    RECT 1.9300 1.7750 3.1950 1.9900 ;
	    RECT 1.5900 1.3200 2.6850 1.5650 ;
	    RECT 1.5900 1.0300 1.7600 1.3200 ;
	    RECT 2.8550 1.1050 3.1950 1.7750 ;
	    RECT 0.0950 0.3200 0.4250 0.8950 ;
	    RECT 1.3850 0.3200 1.7600 1.0300 ;
	    RECT 1.9300 0.8950 3.1950 1.1050 ;
	    RECT 1.9300 0.3200 2.2600 0.8950 ;
   END
END efs8hd_clkdlybuf4s18_1
MACRO efs8hd_clkdlybuf4s18_2
   CLASS CORE ;
   FOREIGN efs8hd_clkdlybuf4s18_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.6800 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 2.7150 1.9050 3.1500 3.0800 ;
	    RECT 2.7150 1.7750 3.1800 1.9050 ;
	    RECT 3.0100 1.1800 3.1800 1.7750 ;
	    RECT 2.9650 0.9750 3.1800 1.1800 ;
	    RECT 2.9650 0.8000 3.1500 0.9750 ;
	    RECT 2.7050 0.3400 3.1500 0.8000 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3450 0.5600 1.6150 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5850 0.1050 0.9150 0.7050 ;
	    RECT 2.1650 0.1050 2.5350 0.7050 ;
	    RECT 3.3200 0.1050 3.5950 0.8050 ;
	    RECT 0.5850 0.0850 3.5950 0.1050 ;
	    RECT 0.0000 -0.0850 3.6800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.6800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.6800 3.4850 ;
	    RECT 0.6000 3.2950 3.5950 3.3150 ;
	    RECT 0.6000 2.2500 0.9300 3.2950 ;
	    RECT 2.1300 2.2500 2.5450 3.2950 ;
	    RECT 3.3200 2.0300 3.5950 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.6800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.0400 0.4300 3.0800 ;
	    RECT 1.1100 2.2500 1.4400 3.0800 ;
	    RECT 0.0850 1.8250 1.0550 2.0400 ;
	    RECT 0.7300 1.1300 1.0550 1.8250 ;
	    RECT 0.0850 0.9200 1.0550 1.1300 ;
	    RECT 1.2700 1.5700 1.4400 2.2500 ;
	    RECT 1.6300 2.0400 1.9600 3.0800 ;
	    RECT 1.6300 1.8250 2.5450 2.0400 ;
	    RECT 1.2700 1.3450 2.2050 1.5700 ;
	    RECT 2.3750 1.5550 2.5450 1.8250 ;
	    RECT 2.3750 1.3450 2.8400 1.5550 ;
	    RECT 0.0850 0.3400 0.4150 0.9200 ;
	    RECT 1.2700 0.7500 1.4400 1.3450 ;
	    RECT 2.3750 1.1300 2.5450 1.3450 ;
	    RECT 1.1600 0.3400 1.4400 0.7500 ;
	    RECT 1.6300 0.9200 2.5450 1.1300 ;
	    RECT 1.6300 0.3400 1.9600 0.9200 ;
   END
END efs8hd_clkdlybuf4s18_2
MACRO efs8hd_clkdlybuf4s25_1
   CLASS CORE ;
   FOREIGN efs8hd_clkdlybuf4s25_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.6800 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 3.0350 1.9550 3.5950 3.0800 ;
	    RECT 3.2300 0.8000 3.5950 1.9550 ;
	    RECT 3.0150 0.3200 3.5950 0.8000 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3450 0.4850 1.6500 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5800 0.1050 0.9100 0.7050 ;
	    RECT 2.2400 0.1050 2.8450 0.7050 ;
	    RECT 0.5800 0.0850 2.8450 0.1050 ;
	    RECT 0.0000 -0.0850 3.6800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.6800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.6800 3.4850 ;
	    RECT 0.6000 3.2950 2.8450 3.3150 ;
	    RECT 0.6000 2.2900 0.9250 3.2950 ;
	    RECT 2.2350 2.2950 2.8450 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.6800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.0750 0.4300 3.0800 ;
	    RECT 1.1950 2.2400 1.6450 3.0800 ;
	    RECT 0.0850 1.8650 1.0050 2.0750 ;
	    RECT 0.6550 1.6200 1.0050 1.8650 ;
	    RECT 0.6550 1.2800 1.1050 1.6200 ;
	    RECT 1.4700 1.5650 1.6450 2.2400 ;
	    RECT 1.8150 2.0800 2.0650 3.0800 ;
	    RECT 1.8150 1.8700 2.7650 2.0800 ;
	    RECT 2.5950 1.6550 2.7650 1.8700 ;
	    RECT 1.4700 1.3450 2.4200 1.5650 ;
	    RECT 0.6550 1.1300 1.0050 1.2800 ;
	    RECT 0.0850 0.9200 1.0050 1.1300 ;
	    RECT 1.4700 1.0700 1.6450 1.3450 ;
	    RECT 2.5950 1.2400 3.0500 1.6550 ;
	    RECT 2.5950 1.1300 2.7650 1.2400 ;
	    RECT 0.0850 0.3200 0.4100 0.9200 ;
	    RECT 1.1750 0.3200 1.6450 1.0700 ;
	    RECT 1.8150 0.9200 2.7650 1.1300 ;
	    RECT 1.8150 0.3200 2.0650 0.9200 ;
   END
END efs8hd_clkdlybuf4s25_1
MACRO efs8hd_clkdlybuf4s25_2
   CLASS CORE ;
   FOREIGN efs8hd_clkdlybuf4s25_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.6800 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 2.7700 2.0300 3.0950 3.0750 ;
	    RECT 2.8650 1.5950 3.0950 2.0300 ;
	    RECT 2.8650 0.9550 3.5950 1.5950 ;
	    RECT 2.8650 0.7700 3.0950 0.9550 ;
	    RECT 2.7700 0.3550 3.0950 0.7700 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.1050 0.4950 2.0200 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5750 0.1050 0.9050 0.5900 ;
	    RECT 2.1350 0.1050 2.4650 0.5800 ;
	    RECT 3.2650 0.1050 3.5950 0.6900 ;
	    RECT 0.5750 0.0850 3.5950 0.1050 ;
	    RECT 0.0000 -0.0850 3.6800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.6800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.6800 3.4850 ;
	    RECT 0.5750 3.2950 3.5950 3.3150 ;
	    RECT 0.5750 2.6550 0.9050 3.2950 ;
	    RECT 2.1350 2.3950 2.4650 3.2950 ;
	    RECT 3.2650 2.0450 3.5950 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.6800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0950 2.4450 0.3450 3.0800 ;
	    RECT 0.0950 2.2300 0.8350 2.4450 ;
	    RECT 0.6650 2.1900 0.8350 2.2300 ;
	    RECT 0.6650 1.6550 1.0050 2.1900 ;
	    RECT 1.1750 1.7800 1.4400 3.0800 ;
	    RECT 1.6950 2.1800 1.9450 3.0800 ;
	    RECT 1.6950 1.8750 2.5950 2.1800 ;
	    RECT 1.2050 1.6550 1.4400 1.7800 ;
	    RECT 0.6650 1.2450 1.0350 1.6550 ;
	    RECT 1.2050 1.2450 2.1650 1.6550 ;
	    RECT 0.6650 0.9350 0.8400 1.2450 ;
	    RECT 1.2050 0.9750 1.4250 1.2450 ;
	    RECT 2.3350 1.0050 2.5950 1.8750 ;
	    RECT 0.0950 0.7650 0.8400 0.9350 ;
	    RECT 0.0950 0.3800 0.3450 0.7650 ;
	    RECT 1.0950 0.3200 1.4250 0.9750 ;
	    RECT 1.6150 0.7950 2.5950 1.0050 ;
	    RECT 1.6150 0.3200 1.9450 0.7950 ;
   END
END efs8hd_clkdlybuf4s25_2
MACRO efs8hd_clkdlybuf4s50_1
   CLASS CORE ;
   FOREIGN efs8hd_clkdlybuf4s50_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.6800 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 3.1900 2.1150 3.5950 3.0800 ;
	    RECT 3.3450 0.8000 3.5950 2.1150 ;
	    RECT 3.1900 0.3200 3.5950 0.8000 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3450 0.5350 1.6150 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5850 0.1050 0.9150 0.7050 ;
	    RECT 2.6900 0.1050 3.0200 0.7500 ;
	    RECT 0.5850 0.0850 3.0200 0.1050 ;
	    RECT 0.0000 -0.0850 3.6800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.6800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.6800 3.4850 ;
	    RECT 0.6000 3.2950 3.0200 3.3150 ;
	    RECT 0.6000 2.2500 0.9300 3.2950 ;
	    RECT 2.6900 2.2950 3.0200 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.6800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.0400 0.4300 3.0800 ;
	    RECT 0.0850 1.8250 1.0550 2.0400 ;
	    RECT 0.7050 1.6450 1.0550 1.8250 ;
	    RECT 1.3800 1.6500 1.7300 3.0800 ;
	    RECT 1.9900 2.0800 2.2400 3.0800 ;
	    RECT 1.9900 1.8700 2.5800 2.0800 ;
	    RECT 2.4100 1.6550 2.5800 1.8700 ;
	    RECT 0.7050 1.2800 1.1350 1.6450 ;
	    RECT 1.3800 1.3400 2.2400 1.6500 ;
	    RECT 0.7050 1.1300 1.0550 1.2800 ;
	    RECT 0.0850 0.9200 1.0550 1.1300 ;
	    RECT 0.0850 0.3200 0.4150 0.9200 ;
	    RECT 1.3800 0.3200 1.7300 1.3400 ;
	    RECT 2.4100 1.2450 3.1750 1.6550 ;
	    RECT 2.4100 1.1250 2.5800 1.2450 ;
	    RECT 1.9900 0.9150 2.5800 1.1250 ;
	    RECT 1.9900 0.3200 2.2400 0.9150 ;
   END
END efs8hd_clkdlybuf4s50_1
MACRO efs8hd_clkdlybuf4s50_2
   CLASS CORE ;
   FOREIGN efs8hd_clkdlybuf4s50_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.1400 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 3.1850 1.9150 3.6250 3.0800 ;
	    RECT 3.3450 0.8000 3.6250 1.9150 ;
	    RECT 3.1850 0.3400 3.6250 0.8000 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3450 0.4800 1.6150 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5850 0.1050 0.9150 0.7050 ;
	    RECT 2.6850 0.1050 3.0150 0.7050 ;
	    RECT 3.7950 0.1050 4.0550 0.7950 ;
	    RECT 0.5850 0.0850 4.0550 0.1050 ;
	    RECT 0.0000 -0.0850 4.1400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.1400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.1400 3.4850 ;
	    RECT 0.6000 3.2950 4.0550 3.3150 ;
	    RECT 0.6000 2.2500 0.9300 3.2950 ;
	    RECT 2.6850 2.2500 3.0150 3.2950 ;
	    RECT 3.7950 2.2500 4.0550 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.1400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.0400 0.4300 3.0800 ;
	    RECT 1.3900 2.2300 1.7950 3.0800 ;
	    RECT 0.0850 1.8200 1.2700 2.0400 ;
	    RECT 0.8500 1.5550 1.2700 1.8200 ;
	    RECT 1.6250 1.5550 1.7950 2.2300 ;
	    RECT 1.9850 2.0400 2.2350 3.0800 ;
	    RECT 1.9850 1.8250 2.6450 2.0400 ;
	    RECT 2.4750 1.6550 2.6450 1.8250 ;
	    RECT 0.7650 1.3450 1.4350 1.5550 ;
	    RECT 1.6250 1.3450 2.3050 1.5550 ;
	    RECT 0.8500 1.1300 1.2700 1.3450 ;
	    RECT 0.0850 0.9200 1.2700 1.1300 ;
	    RECT 1.6250 1.1250 1.7950 1.3450 ;
	    RECT 2.4750 1.2450 3.1750 1.6550 ;
	    RECT 2.4750 1.1300 2.6450 1.2450 ;
	    RECT 0.0850 0.3400 0.4150 0.9200 ;
	    RECT 1.4400 0.3400 1.7950 1.1250 ;
	    RECT 1.9850 0.9200 2.6450 1.1300 ;
	    RECT 1.9850 0.3400 2.2350 0.9200 ;
   END
END efs8hd_clkdlybuf4s50_2
MACRO efs8hd_clkinv_16
   CLASS CORE ;
   FOREIGN efs8hd_clkinv_16 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 11.0400 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.3450 1.1050 2.1550 1.5950 ;
	    RECT 8.9300 1.1200 10.7100 1.5950 ;
         LAYER met1 ;
	    RECT 1.4650 1.5750 2.2150 1.6300 ;
	    RECT 9.2850 1.5750 10.0350 1.6300 ;
	    RECT 1.4650 1.4000 10.0350 1.5750 ;
	    RECT 1.4650 1.3450 2.2150 1.4000 ;
	    RECT 9.2850 1.3450 10.0350 1.4000 ;
      END
   END A
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5750 2.0800 0.8300 3.0800 ;
	    RECT 1.4350 2.0800 1.6900 3.0650 ;
	    RECT 2.3250 2.0800 2.5500 3.0800 ;
	    RECT 3.1550 2.0800 3.4100 3.0650 ;
	    RECT 4.0150 2.0800 4.2550 3.0650 ;
	    RECT 4.9050 2.0800 5.2800 3.0650 ;
	    RECT 5.9250 2.0800 6.1750 3.0650 ;
	    RECT 6.7850 2.0800 7.0350 3.0650 ;
	    RECT 7.6450 2.0800 7.8950 3.0650 ;
	    RECT 8.5050 2.0800 8.7550 3.0650 ;
	    RECT 9.3650 2.0800 9.6050 3.0650 ;
	    RECT 10.2250 2.0800 10.4800 3.0650 ;
	    RECT 0.5750 1.8200 10.4800 2.0800 ;
	    RECT 2.3250 1.7700 8.7550 1.8200 ;
	    RECT 2.3250 0.3500 2.5500 1.7700 ;
	    RECT 3.1550 0.3500 3.4100 1.7700 ;
	    RECT 4.0150 0.3500 4.2550 1.7700 ;
	    RECT 4.9050 0.3500 5.2550 1.7700 ;
	    RECT 5.9250 0.3500 6.1750 1.7700 ;
	    RECT 6.7850 0.3500 7.0350 1.7700 ;
	    RECT 7.6450 0.3500 7.8950 1.7700 ;
	    RECT 8.5050 0.3500 8.7550 1.7700 ;
      END
   END Y
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 1.8550 0.1050 2.1250 0.7650 ;
	    RECT 2.7200 0.1050 2.9850 0.7650 ;
	    RECT 3.5800 0.1050 3.8450 0.7650 ;
	    RECT 4.4650 0.1050 4.7300 0.7650 ;
	    RECT 5.4900 0.1050 5.7550 0.7650 ;
	    RECT 6.3500 0.1050 6.5750 0.7650 ;
	    RECT 7.2100 0.1050 7.4750 0.7650 ;
	    RECT 8.0700 0.1050 8.3350 0.7650 ;
	    RECT 8.9300 0.1050 9.1950 0.7650 ;
	    RECT 1.8550 0.0850 9.1950 0.1050 ;
	    RECT 0.0000 -0.0850 11.0400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 11.0400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 11.0400 3.4850 ;
	    RECT 0.1400 3.2950 10.9100 3.3150 ;
	    RECT 0.1400 1.8700 0.4050 3.2950 ;
	    RECT 1.0000 2.2950 1.2600 3.2950 ;
	    RECT 1.8650 2.2950 2.1200 3.2950 ;
	    RECT 2.7200 2.2950 2.9800 3.2950 ;
	    RECT 3.5850 2.2950 3.8400 3.2950 ;
	    RECT 4.4650 2.2950 4.7200 3.2950 ;
	    RECT 5.4900 2.6500 5.7500 3.2950 ;
	    RECT 5.4900 2.2950 5.7450 2.6500 ;
	    RECT 6.3550 2.2950 6.6100 3.2950 ;
	    RECT 7.2150 2.2950 7.4700 3.2950 ;
	    RECT 8.0750 2.2950 8.3300 3.2950 ;
	    RECT 8.9350 2.2950 9.1900 3.2950 ;
	    RECT 9.7950 2.2950 10.0500 3.2950 ;
	    RECT 10.6500 2.2950 10.9100 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 11.0400 3.7000 ;
      END
   END vpwr
END efs8hd_clkinv_16
MACRO efs8hd_clkinv_1
   CLASS CORE ;
   FOREIGN efs8hd_clkinv_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 1.3800 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.4700 0.3250 1.6550 ;
      END
   END A
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5150 1.6150 0.8450 3.0800 ;
	    RECT 0.5150 0.9500 1.2950 1.6150 ;
	    RECT 0.5150 0.3200 0.8400 0.9500 ;
      END
   END Y
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 1.0100 0.0850 1.2950 0.7400 ;
	    RECT 0.0000 -0.0850 1.3800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 1.3800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 1.3800 3.4850 ;
	    RECT 0.0850 3.2950 1.2950 3.3150 ;
	    RECT 0.0850 2.0800 0.3450 3.2950 ;
	    RECT 1.0150 2.0800 1.2950 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 1.3800 3.7000 ;
      END
   END vpwr
END efs8hd_clkinv_1
MACRO efs8hd_clkinv_2
   CLASS CORE ;
   FOREIGN efs8hd_clkinv_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 1.8400 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.1550 2.0400 0.4100 3.0450 ;
	    RECT 1.0100 2.0400 1.2700 3.0450 ;
	    RECT 0.1550 1.8250 1.7550 2.0400 ;
	    RECT 1.4750 1.1200 1.7550 1.8250 ;
	    RECT 1.0250 0.9050 1.7550 1.1200 ;
	    RECT 1.0250 0.3500 1.2500 0.9050 ;
      END
   END Y
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3300 1.3050 1.6150 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5600 0.1050 0.8550 0.7650 ;
	    RECT 1.4200 0.1050 1.7500 0.6950 ;
	    RECT 0.5600 0.0850 1.7500 0.1050 ;
	    RECT 0.0000 -0.0850 1.8400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 1.8400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 1.8400 3.4850 ;
	    RECT 0.5800 3.2950 1.6950 3.3150 ;
	    RECT 0.5800 2.2500 0.8400 3.2950 ;
	    RECT 1.4400 2.2500 1.6950 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 1.8400 3.7000 ;
      END
   END vpwr
END efs8hd_clkinv_2
MACRO efs8hd_clkinv_4
   CLASS CORE ;
   FOREIGN efs8hd_clkinv_4 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.2200 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.6050 2.0400 0.8600 3.0450 ;
	    RECT 1.4650 2.0400 1.7200 3.0450 ;
	    RECT 2.3200 2.0400 2.5800 3.0450 ;
	    RECT 0.1050 1.8250 3.1350 2.0400 ;
	    RECT 0.1050 1.1200 0.2750 1.8250 ;
	    RECT 2.8350 1.1200 3.1350 1.8250 ;
	    RECT 0.1050 0.9050 3.1350 1.1200 ;
	    RECT 1.0300 0.3500 1.2900 0.9050 ;
	    RECT 1.8900 0.3500 2.1450 0.9050 ;
      END
   END Y
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.4450 1.3300 2.6600 1.6150 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5650 0.1050 0.8600 0.6950 ;
	    RECT 1.4600 0.1050 1.7200 0.6950 ;
	    RECT 2.3150 0.1050 2.6150 0.6950 ;
	    RECT 0.5650 0.0850 2.6150 0.1050 ;
	    RECT 0.0000 -0.0850 3.2200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.2200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.2200 3.4850 ;
	    RECT 0.0850 3.2950 3.1350 3.3150 ;
	    RECT 0.0850 2.2500 0.4300 3.2950 ;
	    RECT 1.0300 2.2500 1.2900 3.2950 ;
	    RECT 1.8900 2.2500 2.1500 3.2950 ;
	    RECT 2.7500 2.2500 3.1350 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.2200 3.7000 ;
      END
   END vpwr
END efs8hd_clkinv_4
MACRO efs8hd_clkinv_8
   CLASS CORE ;
   FOREIGN efs8hd_clkinv_8 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.9800 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5650 2.0400 0.8050 3.0450 ;
	    RECT 1.4050 2.0400 1.6450 3.0450 ;
	    RECT 2.2450 2.0400 2.4950 3.0450 ;
	    RECT 3.0800 2.0400 3.3250 3.0450 ;
	    RECT 3.9200 2.0400 4.1750 3.0450 ;
	    RECT 4.7650 2.0400 5.0050 3.0450 ;
	    RECT 0.1150 1.8250 5.4400 2.0400 ;
	    RECT 0.1150 1.0800 0.2850 1.8250 ;
	    RECT 5.1700 1.0800 5.4400 1.8250 ;
	    RECT 0.1150 0.8700 5.4400 1.0800 ;
	    RECT 1.5350 0.3500 1.7250 0.8700 ;
	    RECT 2.3950 0.3500 2.5850 0.8700 ;
	    RECT 3.2550 0.3500 3.4450 0.8700 ;
	    RECT 4.1150 0.3500 4.3050 0.8700 ;
      END
   END Y
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.4550 1.2950 4.8650 1.6150 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 1.0350 0.1050 1.3650 0.6550 ;
	    RECT 1.8950 0.1050 2.2250 0.6550 ;
	    RECT 2.7550 0.1050 3.0850 0.6550 ;
	    RECT 3.6150 0.1050 3.9450 0.6550 ;
	    RECT 4.4750 0.1050 4.8050 0.6550 ;
	    RECT 1.0350 0.0850 4.8050 0.1050 ;
	    RECT 0.0000 -0.0850 5.9800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.9800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.9800 3.4850 ;
	    RECT 0.1350 3.2950 5.4300 3.3150 ;
	    RECT 0.1350 2.2500 0.3950 3.2950 ;
	    RECT 0.9750 2.2500 1.2350 3.2950 ;
	    RECT 1.8150 2.2500 2.0750 3.2950 ;
	    RECT 2.6650 2.2500 2.9100 3.2950 ;
	    RECT 3.4950 2.2500 3.7500 3.2950 ;
	    RECT 4.3450 2.2500 4.5950 3.2950 ;
	    RECT 5.1750 2.2500 5.4300 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.9800 3.7000 ;
      END
   END vpwr
END efs8hd_clkinv_8
MACRO efs8hd_clkinvlp_2
   CLASS CORE ;
   FOREIGN efs8hd_clkinvlp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 1.8400 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.8100 0.9400 1.2350 3.0700 ;
	    RECT 0.8100 0.3950 1.4450 0.9400 ;
      END
   END Y
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.1450 1.1050 0.6000 2.0800 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.2950 0.0850 0.6250 0.9300 ;
	    RECT 0.0000 -0.0850 1.8400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 1.8400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 1.8400 3.4850 ;
	    RECT 0.2250 3.2800 1.7400 3.3150 ;
	    RECT 0.2250 2.2950 0.5550 3.2800 ;
	    RECT 1.4400 1.8200 1.7400 3.2800 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 1.8400 3.7000 ;
      END
   END vpwr
END efs8hd_clkinvlp_2
MACRO efs8hd_clkinvlp_4
   CLASS CORE ;
   FOREIGN efs8hd_clkinvlp_4 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 2.7600 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5950 1.6200 0.9550 3.0800 ;
	    RECT 1.6850 1.6200 2.0150 3.0800 ;
	    RECT 0.5950 1.2700 2.0150 1.6200 ;
	    RECT 0.5950 0.8500 0.9550 1.2700 ;
	    RECT 0.5950 0.3200 1.2150 0.8500 ;
      END
   END Y
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.7650 0.4250 1.6550 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0950 0.1050 0.4250 0.5950 ;
	    RECT 1.6750 0.1050 2.0050 0.9700 ;
	    RECT 0.0950 0.0850 2.0050 0.1050 ;
	    RECT 0.0000 -0.0850 2.7600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 2.7600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 2.7600 3.4850 ;
	    RECT 0.0950 3.2950 2.5450 3.3150 ;
	    RECT 0.0950 1.8700 0.4250 3.2950 ;
	    RECT 1.1550 1.8300 1.4850 3.2950 ;
	    RECT 2.2150 1.8300 2.5450 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 2.7600 3.7000 ;
      END
   END vpwr
END efs8hd_clkinvlp_4
MACRO efs8hd_conb_1
   CLASS CORE ;
   FOREIGN efs8hd_conb_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 1.3800 BY 3.4000 ;
   SITE unitehd ;
   PIN HI
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 1.3800 3.4850 ;
	    RECT 0.2750 2.3850 0.6050 3.3150 ;
	    RECT 0.0850 0.3150 0.6050 2.1750 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 1.3800 3.7000 ;
      END
   END HI
   PIN LO
      PORT
         LAYER li1 ;
	    RECT 0.7750 1.1400 1.2950 3.0800 ;
	    RECT 0.7750 0.0850 1.1150 0.9300 ;
	    RECT 0.0000 -0.0850 1.3800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 1.3800 0.3000 ;
      END
   END LO
END efs8hd_conb_1
MACRO efs8hd_decap_12
   CLASS CORE ;
   FOREIGN efs8hd_decap_12 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.5200 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.0650 2.6650 1.7150 ;
	    RECT 0.0850 0.0850 5.4300 1.0650 ;
	    RECT 0.0000 -0.0850 5.5200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.5200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.5200 3.4850 ;
	    RECT 0.0850 1.9300 5.4300 3.3150 ;
	    RECT 2.8350 1.2800 5.4300 1.9300 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.5200 3.7000 ;
      END
   END vpwr
END efs8hd_decap_12
MACRO efs8hd_decap_3
   CLASS CORE ;
   FOREIGN efs8hd_decap_3 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 1.3800 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.0400 0.6050 1.7150 ;
	    RECT 0.0850 0.0850 1.2950 1.0400 ;
	    RECT 0.0000 -0.0850 1.3800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 1.3800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 1.3800 3.4850 ;
	    RECT 0.0850 1.9300 1.2950 3.3150 ;
	    RECT 0.7750 1.2550 1.2950 1.9300 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 1.3800 3.7000 ;
      END
   END vpwr
END efs8hd_decap_3
MACRO efs8hd_decap_4
   CLASS CORE ;
   FOREIGN efs8hd_decap_4 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 1.8400 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.0650 0.8350 1.7150 ;
	    RECT 0.0850 0.0850 1.7550 1.0650 ;
	    RECT 0.0000 -0.0850 1.8400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 1.8400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 1.8400 3.4850 ;
	    RECT 0.0850 1.9300 1.7550 3.3150 ;
	    RECT 1.0050 1.2800 1.7550 1.9300 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 1.8400 3.7000 ;
      END
   END vpwr
END efs8hd_decap_4
MACRO efs8hd_decap_6
   CLASS CORE ;
   FOREIGN efs8hd_decap_6 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 2.7600 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.0650 1.2950 1.7150 ;
	    RECT 0.0850 0.0850 2.6750 1.0650 ;
	    RECT 0.0000 -0.0850 2.7600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 2.7600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 2.7600 3.4850 ;
	    RECT 0.0850 1.9300 2.6750 3.3150 ;
	    RECT 1.4650 1.2800 2.6750 1.9300 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 2.7600 3.7000 ;
      END
   END vpwr
END efs8hd_decap_6
MACRO efs8hd_decap_8
   CLASS CORE ;
   FOREIGN efs8hd_decap_8 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.6800 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.0650 1.7350 1.7150 ;
	    RECT 0.0850 0.0850 3.5950 1.0650 ;
	    RECT 0.0000 -0.0850 3.6800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.6800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.6800 3.4850 ;
	    RECT 0.0850 1.9300 3.5950 3.3150 ;
	    RECT 1.9050 1.2800 3.5950 1.9300 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.6800 3.7000 ;
      END
   END vpwr
END efs8hd_decap_8
MACRO efs8hd_dfbbn_2
   CLASS CORE ;
   FOREIGN efs8hd_dfbbn_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 12.8800 BY 3.4000 ;
   SITE unitehd ;
   PIN RESETB
      PORT
         LAYER li1 ;
	    RECT 9.2500 1.3700 9.7300 1.6550 ;
      END
   END RESETB
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.4450 0.1050 1.7850 0.5800 ;
	    RECT 3.5800 0.1050 3.7500 0.6550 ;
	    RECT 5.3600 0.1050 5.6900 0.5800 ;
	    RECT 7.2750 0.1050 7.5350 0.6550 ;
	    RECT 9.7400 0.1050 10.0700 1.0050 ;
	    RECT 10.6800 0.1050 10.9100 1.1050 ;
	    RECT 11.6500 0.1050 11.9450 0.6800 ;
	    RECT 12.5150 0.1050 12.7950 1.1050 ;
	    RECT 0.0000 -0.1050 12.8800 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 12.8800 0.3000 ;
      END
   END vgnd
   PIN CLKN
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.2200 0.4400 2.0300 ;
      END
   END CLKN
   PIN SETB
      PORT
         LAYER li1 ;
	    RECT 3.6000 1.2050 3.9300 1.3300 ;
	    RECT 3.6000 0.9200 4.0100 1.2050 ;
	    RECT 7.4700 0.9200 7.8450 1.3300 ;
         LAYER met1 ;
	    RECT 3.7800 1.1500 4.0700 1.2050 ;
	    RECT 7.4600 1.1500 7.7500 1.2050 ;
	    RECT 3.7800 0.9750 7.7500 1.1500 ;
	    RECT 3.7800 0.9200 4.0700 0.9750 ;
	    RECT 7.4600 0.9200 7.7500 0.9750 ;
      END
   END SETB
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 12.1150 1.8050 12.3450 3.0800 ;
	    RECT 12.1600 1.0300 12.3450 1.8050 ;
	    RECT 12.1150 0.3200 12.3450 1.0300 ;
      END
   END Q
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 12.8800 3.5050 ;
	    RECT 0.5150 2.6700 0.8450 3.2950 ;
	    RECT 1.4450 2.6700 1.7850 3.2950 ;
	    RECT 3.4200 2.7550 3.8000 3.2950 ;
	    RECT 4.8900 2.3950 5.2200 3.2950 ;
	    RECT 7.3350 2.8200 7.7150 3.2950 ;
	    RECT 8.6550 2.8200 10.0700 3.2950 ;
	    RECT 10.6800 1.8300 10.9100 3.2950 ;
	    RECT 11.6500 2.2050 11.9450 3.2950 ;
	    RECT 12.5150 1.8300 12.7950 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 12.8800 3.7000 ;
      END
   END vpwr
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.7600 1.2550 2.1700 2.0300 ;
      END
   END D
   PIN QN
      PORT
         LAYER li1 ;
	    RECT 10.2400 2.0400 10.5000 3.0800 ;
	    RECT 10.3200 0.8950 10.5000 2.0400 ;
	    RECT 10.2400 0.3200 10.5000 0.8950 ;
      END
   END QN
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.4550 0.3450 3.0800 ;
	    RECT 0.0850 2.2450 0.8400 2.4550 ;
	    RECT 0.6100 1.0050 0.8400 2.2450 ;
	    RECT 0.0850 0.7950 0.8400 1.0050 ;
	    RECT 0.0850 0.4300 0.3450 0.7950 ;
	    RECT 1.0150 0.4300 1.2400 3.0800 ;
	    RECT 1.9550 2.4550 2.1250 3.0800 ;
	    RECT 2.3500 2.8150 3.1800 3.0250 ;
	    RECT 1.4200 2.2450 2.1250 2.4550 ;
	    RECT 1.4200 1.0300 1.5900 2.2450 ;
	    RECT 2.3400 1.9700 2.8400 2.4450 ;
	    RECT 1.4200 0.7950 2.1250 1.0300 ;
	    RECT 2.3400 0.8800 2.5600 1.9700 ;
	    RECT 3.0100 1.7550 3.1800 2.8150 ;
	    RECT 4.1000 2.5450 4.2700 2.9700 ;
	    RECT 6.2650 2.8150 7.0950 3.0250 ;
	    RECT 3.3500 2.2300 4.7000 2.5450 ;
	    RECT 3.3500 1.9700 3.6000 2.2300 ;
	    RECT 4.1100 1.7550 4.3600 1.8550 ;
	    RECT 3.0100 1.5450 4.3600 1.7550 ;
	    RECT 3.0100 1.4950 3.4100 1.5450 ;
	    RECT 2.7400 0.8050 3.0700 1.2700 ;
	    RECT 1.9550 0.3800 2.1250 0.7950 ;
	    RECT 3.2400 0.5800 3.4100 1.4950 ;
	    RECT 4.1400 1.4450 4.3600 1.5450 ;
	    RECT 4.5300 1.3300 4.7000 2.2300 ;
	    RECT 4.8700 1.7700 5.8750 2.0700 ;
	    RECT 6.0750 1.9700 6.3100 2.4800 ;
	    RECT 4.8700 1.5450 5.2000 1.7700 ;
	    RECT 6.5500 1.6300 6.7550 2.3800 ;
	    RECT 5.5100 1.3300 5.8400 1.5450 ;
	    RECT 4.5300 1.1200 5.8400 1.3300 ;
	    RECT 6.1350 1.4050 6.7550 1.6300 ;
	    RECT 6.9250 1.7550 7.0950 2.8150 ;
	    RECT 7.9550 2.6050 8.1250 2.9700 ;
	    RECT 7.2650 2.3950 10.0700 2.6050 ;
	    RECT 7.2650 1.9700 7.5150 2.3950 ;
	    RECT 6.9250 1.5450 8.2750 1.7550 ;
	    RECT 4.5300 0.9550 4.7500 1.1200 ;
	    RECT 4.4200 0.7450 4.7500 0.9550 ;
	    RECT 2.4150 0.3300 3.4100 0.5800 ;
	    RECT 3.9200 0.5300 4.2500 0.6800 ;
	    RECT 4.9200 0.5300 5.1700 0.8950 ;
	    RECT 6.1350 0.8800 6.4200 1.4050 ;
	    RECT 6.9250 0.5800 7.0950 1.5450 ;
	    RECT 8.0550 1.3450 8.2750 1.5450 ;
	    RECT 8.4450 0.9750 8.6250 2.3950 ;
	    RECT 8.2950 0.7450 8.6250 0.9750 ;
	    RECT 8.7950 1.9700 9.5700 2.1800 ;
	    RECT 8.7950 1.1550 9.0700 1.9700 ;
	    RECT 9.9000 1.6550 10.0700 2.3950 ;
	    RECT 11.2150 1.6550 11.4700 3.0200 ;
	    RECT 9.9000 1.2450 10.1400 1.6550 ;
	    RECT 11.2150 1.2450 11.9900 1.6550 ;
	    RECT 8.7950 0.9450 9.5000 1.1550 ;
	    RECT 3.9200 0.3200 5.1700 0.5300 ;
	    RECT 6.3300 0.3300 7.0950 0.5800 ;
	    RECT 7.7950 0.5300 8.1250 0.6800 ;
	    RECT 8.7950 0.5300 8.9650 0.7300 ;
	    RECT 7.7950 0.3200 8.9650 0.5300 ;
	    RECT 9.2800 0.3300 9.5000 0.9450 ;
	    RECT 11.2150 0.3200 11.4700 1.2450 ;
         LAYER met1 ;
	    RECT 1.0100 2.4250 1.3000 2.4800 ;
	    RECT 2.4000 2.4250 2.6900 2.4800 ;
	    RECT 6.0800 2.4250 6.3700 2.4800 ;
	    RECT 1.0100 2.2500 6.3700 2.4250 ;
	    RECT 1.0100 2.1950 1.3000 2.2500 ;
	    RECT 2.4000 2.1950 2.6900 2.2500 ;
	    RECT 6.0800 2.1950 6.3700 2.2500 ;
	    RECT 5.6200 2.0000 5.9100 2.0550 ;
	    RECT 8.8400 2.0000 9.1300 2.0550 ;
	    RECT 5.6200 1.8250 9.1300 2.0000 ;
	    RECT 5.6200 1.7700 5.9100 1.8250 ;
	    RECT 8.8400 1.7700 9.1300 1.8250 ;
	    RECT 6.0800 1.5750 6.3700 1.6300 ;
	    RECT 2.9350 1.4000 6.3700 1.5750 ;
	    RECT 2.9350 1.2050 3.1300 1.4000 ;
	    RECT 6.0800 1.3450 6.3700 1.4000 ;
	    RECT 0.5500 1.1500 0.8400 1.2050 ;
	    RECT 2.8400 1.1500 3.1300 1.2050 ;
	    RECT 0.5500 0.9750 3.1300 1.1500 ;
	    RECT 0.5500 0.9200 0.8400 0.9750 ;
	    RECT 2.8400 0.9200 3.1300 0.9750 ;
   END
END efs8hd_dfbbn_2
MACRO efs8hd_dfrbp_2
   CLASS CORE ;
   FOREIGN efs8hd_dfrbp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 11.0400 BY 3.4000 ;
   SITE unitehd ;
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 9.1600 0.3300 9.4950 2.1200 ;
      END
   END Q
   PIN QN
      PORT
         LAYER li1 ;
	    RECT 10.1200 2.6000 10.4200 3.0800 ;
	    RECT 10.0300 1.9200 10.4200 2.6000 ;
	    RECT 10.2500 1.0300 10.4200 1.9200 ;
	    RECT 10.0400 0.3900 10.4200 1.0300 ;
      END
   END QN
   PIN RESETB
      PORT
         LAYER li1 ;
	    RECT 7.1050 1.2950 7.6450 1.7550 ;
	    RECT 3.8050 0.9550 4.5950 1.2700 ;
	    RECT 7.4050 0.7950 7.6450 1.2950 ;
         LAYER met1 ;
	    RECT 7.0450 1.2050 7.3350 1.6000 ;
	    RECT 3.7450 1.1500 4.3950 1.2050 ;
	    RECT 7.0450 1.1500 7.6350 1.2050 ;
	    RECT 3.7450 0.9750 7.6350 1.1500 ;
	    RECT 3.7450 0.9200 4.3950 0.9750 ;
	    RECT 7.3450 0.9200 7.6350 0.9750 ;
      END
   END RESETB
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.3550 2.0800 1.6800 3.0650 ;
	    RECT 1.4150 0.7700 1.8750 2.0800 ;
      END
   END D
   PIN CLK
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.2200 0.4400 2.0300 ;
      END
   END CLK
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.5450 0.1050 1.8750 0.5550 ;
	    RECT 4.4750 0.1050 4.8050 0.6800 ;
	    RECT 6.7050 0.1050 6.8950 0.6550 ;
	    RECT 8.7550 0.1050 8.9900 0.6800 ;
	    RECT 9.7000 0.1050 9.8700 1.0300 ;
	    RECT 10.5900 0.1050 10.7600 1.1650 ;
	    RECT 0.0000 -0.1050 11.0400 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 11.0400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 11.0400 3.5050 ;
	    RECT 0.5150 2.6700 0.8450 3.2950 ;
	    RECT 1.8500 2.7200 2.1000 3.2950 ;
	    RECT 3.9900 2.7550 4.3200 3.2950 ;
	    RECT 4.9550 2.7200 5.3250 3.2950 ;
	    RECT 6.9400 2.7200 7.1900 3.2950 ;
	    RECT 7.7100 2.8200 8.0550 3.2950 ;
	    RECT 8.7300 2.7550 9.0700 3.2950 ;
	    RECT 9.6200 2.8200 9.9500 3.2950 ;
	    RECT 10.5900 1.8050 10.7600 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 11.0400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0900 2.4550 0.3450 3.0800 ;
	    RECT 0.0900 2.2450 0.8400 2.4550 ;
	    RECT 0.6100 1.0050 0.8400 2.2450 ;
	    RECT 0.0900 0.7950 0.8400 1.0050 ;
	    RECT 0.0900 0.4300 0.3450 0.7950 ;
	    RECT 1.0150 0.4300 1.1850 3.0800 ;
	    RECT 2.2700 2.6700 2.5200 3.0800 ;
	    RECT 2.7350 2.6700 3.4150 3.0800 ;
	    RECT 2.2700 2.5050 2.4400 2.6700 ;
	    RECT 2.0450 2.2950 2.4400 2.5050 ;
	    RECT 2.0450 0.5950 2.2150 2.2950 ;
	    RECT 2.6100 1.9700 3.0750 2.4550 ;
	    RECT 2.3850 0.9550 2.7350 1.7300 ;
	    RECT 2.9050 1.2300 3.0750 1.9700 ;
	    RECT 3.2450 1.6950 3.4150 2.6700 ;
	    RECT 3.5850 2.5450 3.7550 2.9700 ;
	    RECT 4.4900 2.5450 4.6600 2.9700 ;
	    RECT 3.5850 2.3300 4.6600 2.5450 ;
	    RECT 5.4950 2.5050 5.6650 3.0800 ;
	    RECT 5.9000 2.6550 6.7700 3.0800 ;
	    RECT 5.1050 2.2950 5.6650 2.5050 ;
	    RECT 5.1050 2.1200 5.2750 2.2950 ;
	    RECT 3.7750 1.9050 5.2750 2.1200 ;
	    RECT 5.9700 2.0800 6.4300 2.4450 ;
	    RECT 3.2450 1.4800 4.9350 1.6950 ;
	    RECT 2.9050 0.9550 3.2600 1.2300 ;
	    RECT 3.4300 0.5950 3.6000 1.4800 ;
	    RECT 4.7650 1.2550 4.9350 1.4800 ;
	    RECT 5.1050 1.0450 5.2750 1.9050 ;
	    RECT 2.0450 0.3800 2.5400 0.5950 ;
	    RECT 2.7450 0.3800 3.6000 0.5950 ;
	    RECT 5.0150 0.5550 5.2750 1.0450 ;
	    RECT 5.4650 2.0700 6.4300 2.0800 ;
	    RECT 6.6000 2.1800 6.7700 2.6550 ;
	    RECT 7.3600 2.6050 7.5300 2.9700 ;
	    RECT 7.3600 2.3950 8.1600 2.6050 ;
	    RECT 5.4650 1.8700 6.1400 2.0700 ;
	    RECT 6.6000 1.9700 7.8200 2.1800 ;
	    RECT 5.4650 0.8800 5.6750 1.8700 ;
	    RECT 6.6000 1.8550 6.7700 1.9700 ;
	    RECT 5.8450 0.8800 6.1950 1.6550 ;
	    RECT 6.3650 1.6450 6.7700 1.8550 ;
	    RECT 7.9900 1.6550 8.1600 2.3950 ;
	    RECT 8.3350 2.5450 8.5600 3.0800 ;
	    RECT 8.3350 2.3300 9.8350 2.5450 ;
	    RECT 8.3350 2.2450 8.9900 2.3300 ;
	    RECT 6.3650 0.6700 6.5350 1.6450 ;
	    RECT 7.9900 1.6200 8.6500 1.6550 ;
	    RECT 6.7050 1.0800 6.9250 1.4300 ;
	    RECT 7.8150 1.3450 8.6500 1.6200 ;
	    RECT 7.8150 1.2450 8.1600 1.3450 ;
	    RECT 6.7050 0.8700 7.2350 1.0800 ;
	    RECT 5.0150 0.3450 5.3650 0.5550 ;
	    RECT 5.5850 0.3200 6.5350 0.6700 ;
	    RECT 7.0650 0.5800 7.2350 0.8700 ;
	    RECT 7.8150 0.5800 7.9850 1.2450 ;
	    RECT 8.8200 1.1050 8.9900 2.2450 ;
	    RECT 9.6650 1.6550 9.8350 2.3300 ;
	    RECT 9.6650 1.2450 10.0800 1.6550 ;
	    RECT 7.0650 0.3700 7.9850 0.5800 ;
	    RECT 8.3350 0.8950 8.9900 1.1050 ;
	    RECT 8.3350 0.4300 8.5850 0.8950 ;
         LAYER met1 ;
	    RECT 0.9550 2.4250 1.2450 2.4800 ;
	    RECT 2.8450 2.4250 3.1350 2.4800 ;
	    RECT 5.9650 2.4250 6.2550 2.4800 ;
	    RECT 0.9550 2.2500 6.2550 2.4250 ;
	    RECT 0.9550 2.1950 1.2450 2.2500 ;
	    RECT 2.8450 2.1950 3.1350 2.2500 ;
	    RECT 5.9650 2.1950 6.2550 2.2500 ;
	    RECT 0.5500 1.5750 0.8400 1.6300 ;
	    RECT 2.3850 1.5750 2.6750 1.6300 ;
	    RECT 5.9650 1.5750 6.2550 1.6300 ;
	    RECT 0.5500 1.4000 6.2550 1.5750 ;
	    RECT 0.5500 1.3450 0.8400 1.4000 ;
	    RECT 2.3850 1.3450 2.6750 1.4000 ;
	    RECT 5.9650 1.3450 6.2550 1.4000 ;
   END
END efs8hd_dfrbp_2
MACRO efs8hd_dfrtp_2
   CLASS CORE ;
   FOREIGN efs8hd_dfrtp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 9.6600 BY 3.4000 ;
   SITE unitehd ;
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 8.8550 1.8050 9.1050 2.9050 ;
	    RECT 8.9000 0.9950 9.1050 1.8050 ;
	    RECT 8.8550 0.3300 9.1050 0.9950 ;
      END
   END Q
   PIN RESETB
      PORT
         LAYER li1 ;
	    RECT 7.1050 1.2950 7.6450 1.7550 ;
	    RECT 3.8050 0.9550 4.5950 1.2700 ;
	    RECT 7.4050 0.7950 7.6450 1.2950 ;
         LAYER met1 ;
	    RECT 7.0450 1.2050 7.3350 1.6000 ;
	    RECT 3.7450 1.1500 4.3950 1.2050 ;
	    RECT 7.0450 1.1500 7.6350 1.2050 ;
	    RECT 3.7450 0.9750 7.6350 1.1500 ;
	    RECT 3.7450 0.9200 4.3950 0.9750 ;
	    RECT 7.3450 0.9200 7.6350 0.9750 ;
      END
   END RESETB
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.3550 2.0800 1.6800 3.0650 ;
	    RECT 1.4150 0.7700 1.8750 2.0800 ;
      END
   END D
   PIN CLK
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.2200 0.4400 2.0300 ;
      END
   END CLK
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.5450 0.1050 1.8750 0.5550 ;
	    RECT 4.4750 0.1050 4.8050 0.6800 ;
	    RECT 6.7050 0.1050 6.8950 0.6550 ;
	    RECT 8.3800 0.1050 8.6850 0.6800 ;
	    RECT 9.2750 0.1050 9.5250 1.0500 ;
	    RECT 0.0000 -0.1050 9.6600 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 9.6600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 9.6600 3.5050 ;
	    RECT 0.5150 2.6700 0.8450 3.2950 ;
	    RECT 1.8500 2.7200 2.1000 3.2950 ;
	    RECT 3.9900 2.7550 4.3200 3.2950 ;
	    RECT 4.9550 2.7200 5.3250 3.2950 ;
	    RECT 6.9400 2.7200 7.1900 3.2950 ;
	    RECT 7.7100 2.8200 8.0400 3.2950 ;
	    RECT 8.3800 1.8700 8.6850 3.2950 ;
	    RECT 9.2750 1.8700 9.5250 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 9.6600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0900 2.4550 0.3450 3.0800 ;
	    RECT 0.0900 2.2450 0.8400 2.4550 ;
	    RECT 0.6100 1.0050 0.8400 2.2450 ;
	    RECT 0.0900 0.7950 0.8400 1.0050 ;
	    RECT 0.0900 0.4300 0.3450 0.7950 ;
	    RECT 1.0150 0.4300 1.1850 3.0800 ;
	    RECT 2.2700 2.6700 2.5200 3.0800 ;
	    RECT 2.7350 2.6700 3.4150 3.0800 ;
	    RECT 2.2700 2.5050 2.4400 2.6700 ;
	    RECT 2.0450 2.2950 2.4400 2.5050 ;
	    RECT 2.0450 0.5950 2.2150 2.2950 ;
	    RECT 2.6100 1.9700 3.0750 2.4550 ;
	    RECT 2.3850 0.9550 2.7350 1.7300 ;
	    RECT 2.9050 1.2300 3.0750 1.9700 ;
	    RECT 3.2450 1.6950 3.4150 2.6700 ;
	    RECT 3.5850 2.5450 3.7550 2.9700 ;
	    RECT 4.4900 2.5450 4.6600 2.9700 ;
	    RECT 3.5850 2.3300 4.6600 2.5450 ;
	    RECT 5.4950 2.5050 5.6650 3.0800 ;
	    RECT 5.9000 2.6550 6.7700 3.0800 ;
	    RECT 5.1050 2.2950 5.6650 2.5050 ;
	    RECT 5.1050 2.1200 5.2750 2.2950 ;
	    RECT 3.7750 1.9050 5.2750 2.1200 ;
	    RECT 5.9700 2.0800 6.4300 2.4450 ;
	    RECT 3.2450 1.4800 4.9350 1.6950 ;
	    RECT 2.9050 0.9550 3.2600 1.2300 ;
	    RECT 3.4300 0.5950 3.6000 1.4800 ;
	    RECT 4.7650 1.2550 4.9350 1.4800 ;
	    RECT 5.1050 1.0450 5.2750 1.9050 ;
	    RECT 2.0450 0.3800 2.5400 0.5950 ;
	    RECT 2.7450 0.3800 3.6000 0.5950 ;
	    RECT 5.0150 0.5550 5.2750 1.0450 ;
	    RECT 5.4650 2.0700 6.4300 2.0800 ;
	    RECT 6.6000 2.1800 6.7700 2.6550 ;
	    RECT 7.3600 2.6050 7.5300 2.9700 ;
	    RECT 7.3600 2.3950 8.1600 2.6050 ;
	    RECT 5.4650 1.8700 6.1400 2.0700 ;
	    RECT 6.6000 1.9700 7.8200 2.1800 ;
	    RECT 5.4650 0.8800 5.6750 1.8700 ;
	    RECT 6.6000 1.8550 6.7700 1.9700 ;
	    RECT 5.8450 0.8800 6.1950 1.6550 ;
	    RECT 6.3650 1.6450 6.7700 1.8550 ;
	    RECT 7.9900 1.6550 8.1600 2.3950 ;
	    RECT 6.3650 0.6700 6.5350 1.6450 ;
	    RECT 7.9900 1.6200 8.7300 1.6550 ;
	    RECT 6.7050 1.0800 6.9250 1.4300 ;
	    RECT 7.8150 1.2450 8.7300 1.6200 ;
	    RECT 6.7050 0.8700 7.2350 1.0800 ;
	    RECT 5.0150 0.3450 5.3650 0.5550 ;
	    RECT 5.5850 0.3200 6.5350 0.6700 ;
	    RECT 7.0650 0.5800 7.2350 0.8700 ;
	    RECT 7.8150 1.0250 8.1400 1.2450 ;
	    RECT 7.8150 0.5800 8.1350 1.0250 ;
	    RECT 7.0650 0.3700 8.1350 0.5800 ;
         LAYER met1 ;
	    RECT 0.9550 2.4250 1.2450 2.4800 ;
	    RECT 2.8450 2.4250 3.1350 2.4800 ;
	    RECT 5.9650 2.4250 6.2550 2.4800 ;
	    RECT 0.9550 2.2500 6.2550 2.4250 ;
	    RECT 0.9550 2.1950 1.2450 2.2500 ;
	    RECT 2.8450 2.1950 3.1350 2.2500 ;
	    RECT 5.9650 2.1950 6.2550 2.2500 ;
	    RECT 0.5500 1.5750 0.8400 1.6300 ;
	    RECT 2.3850 1.5750 2.6750 1.6300 ;
	    RECT 5.9650 1.5750 6.2550 1.6300 ;
	    RECT 0.5500 1.4000 6.2550 1.5750 ;
	    RECT 0.5500 1.3450 0.8400 1.4000 ;
	    RECT 2.3850 1.3450 2.6750 1.4000 ;
	    RECT 5.9650 1.3450 6.2550 1.4000 ;
   END
END efs8hd_dfrtp_2
MACRO efs8hd_dfsbp_2
   CLASS CORE ;
   FOREIGN efs8hd_dfsbp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 11.0400 BY 3.4000 ;
   SITE unitehd ;
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 10.1500 2.0800 10.4800 3.0800 ;
	    RECT 10.1500 1.8700 10.9150 2.0800 ;
	    RECT 10.3600 1.0550 10.9150 1.8700 ;
	    RECT 10.3450 1.0300 10.9150 1.0550 ;
	    RECT 10.2300 0.9000 10.9150 1.0300 ;
	    RECT 10.2300 0.3200 10.4800 0.9000 ;
      END
   END Q
   PIN QN
      PORT
         LAYER li1 ;
	    RECT 8.3700 0.3200 8.7000 3.0800 ;
      END
   END QN
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.7700 1.2550 2.1800 2.0300 ;
      END
   END D
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 11.0400 3.5050 ;
	    RECT 0.5150 2.6700 0.8450 3.2950 ;
	    RECT 1.4550 2.6700 1.7850 3.2950 ;
	    RECT 3.4300 2.8200 3.8100 3.2950 ;
	    RECT 4.3300 2.8200 4.6600 3.2950 ;
	    RECT 5.9300 2.8200 6.3400 3.2950 ;
	    RECT 7.0100 2.4300 7.3400 3.2950 ;
	    RECT 8.0200 1.8500 8.2000 3.2950 ;
	    RECT 8.8700 1.8500 9.1200 3.2950 ;
	    RECT 9.8100 1.8700 9.9800 3.2950 ;
	    RECT 10.6500 2.2950 10.9150 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 11.0400 3.7000 ;
      END
   END vpwr
   PIN SETB
      PORT
         LAYER li1 ;
	    RECT 3.6100 0.9200 4.0200 1.3300 ;
	    RECT 6.6600 1.2550 6.9900 1.3300 ;
	    RECT 6.6600 0.9200 7.3200 1.2550 ;
         LAYER met1 ;
	    RECT 3.7650 1.1500 4.0550 1.2050 ;
	    RECT 6.9850 1.1500 7.2750 1.2050 ;
	    RECT 3.7650 0.9750 7.2750 1.1500 ;
	    RECT 3.7650 0.9200 4.0550 0.9750 ;
	    RECT 6.9850 0.9200 7.2750 0.9750 ;
      END
   END SETB
   PIN CLK
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.2200 0.4400 2.0300 ;
      END
   END CLK
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.4550 0.1050 1.7850 0.5800 ;
	    RECT 3.6100 0.1050 4.0200 0.6550 ;
	    RECT 4.7400 0.1050 5.0800 0.6800 ;
	    RECT 6.6700 0.1050 7.3300 0.7050 ;
	    RECT 8.0200 0.1050 8.2000 1.1300 ;
	    RECT 8.8700 0.1050 9.1200 1.1300 ;
	    RECT 9.7300 0.1050 10.0600 1.0300 ;
	    RECT 10.6500 0.1050 10.9150 0.6900 ;
	    RECT 0.0000 -0.1050 11.0400 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 11.0400 0.3000 ;
      END
   END vgnd
   OBS
         LAYER li1 ;
	    RECT 0.1750 2.4550 0.3450 3.0800 ;
	    RECT 0.1750 2.2450 0.8400 2.4550 ;
	    RECT 0.6100 1.0050 0.8400 2.2450 ;
	    RECT 0.1750 0.7950 0.8400 1.0050 ;
	    RECT 0.1750 0.4300 0.3450 0.7950 ;
	    RECT 1.0150 0.4300 1.2400 3.0800 ;
	    RECT 1.9550 2.4550 2.1250 3.0800 ;
	    RECT 2.3600 2.8150 3.1900 3.0250 ;
	    RECT 1.4300 2.2450 2.1250 2.4550 ;
	    RECT 1.4300 1.0300 1.6000 2.2450 ;
	    RECT 2.3500 1.9700 2.8500 2.4450 ;
	    RECT 1.4300 0.7950 2.1250 1.0300 ;
	    RECT 2.3500 0.8800 2.5700 1.9700 ;
	    RECT 3.0200 1.7550 3.1900 2.8150 ;
	    RECT 3.9900 2.6050 4.1600 2.9700 ;
	    RECT 5.1100 2.7050 5.7600 3.0200 ;
	    RECT 5.5900 2.6050 5.7600 2.7050 ;
	    RECT 6.5400 2.6050 6.7800 2.9700 ;
	    RECT 3.3600 2.2950 4.7100 2.6050 ;
	    RECT 3.3600 1.9700 3.6100 2.2950 ;
	    RECT 4.1200 1.7550 4.3700 1.9550 ;
	    RECT 3.0200 1.5450 4.3700 1.7550 ;
	    RECT 3.0200 1.4950 3.4400 1.5450 ;
	    RECT 2.7500 0.8050 3.1000 1.2700 ;
	    RECT 1.9550 0.3800 2.1250 0.7950 ;
	    RECT 3.2700 0.5800 3.4400 1.4950 ;
	    RECT 4.5400 1.3300 4.7100 2.2950 ;
	    RECT 2.4250 0.3300 3.4400 0.5800 ;
	    RECT 4.3100 0.9050 4.7100 1.3300 ;
	    RECT 4.9000 2.0700 5.4000 2.4550 ;
	    RECT 5.5900 2.3950 6.7800 2.6050 ;
	    RECT 4.9000 1.1200 5.0700 2.0700 ;
	    RECT 5.2400 1.3300 5.4200 1.8450 ;
	    RECT 5.5900 1.7550 5.7600 2.3950 ;
	    RECT 7.5100 2.2050 7.6800 2.9700 ;
	    RECT 7.5100 2.1800 7.8300 2.2050 ;
	    RECT 5.9300 1.9700 7.8300 2.1800 ;
	    RECT 5.5900 1.5450 7.4700 1.7550 ;
	    RECT 5.8200 1.1200 6.1500 1.2700 ;
	    RECT 4.9000 0.9050 6.1500 1.1200 ;
	    RECT 4.3100 0.3700 4.5600 0.9050 ;
	    RECT 6.3200 0.5950 6.4900 1.5450 ;
	    RECT 7.1400 1.4700 7.4700 1.5450 ;
	    RECT 7.6400 0.8500 7.8300 1.9700 ;
	    RECT 5.6400 0.3800 6.4900 0.5950 ;
	    RECT 7.5100 0.4400 7.8300 0.8500 ;
	    RECT 9.3100 1.6550 9.6400 3.0800 ;
	    RECT 9.3100 1.2450 10.1900 1.6550 ;
	    RECT 9.3100 0.3200 9.5600 1.2450 ;
         LAYER met1 ;
	    RECT 0.5850 2.4250 0.8750 2.4800 ;
	    RECT 2.3850 2.4250 2.6750 2.4800 ;
	    RECT 5.1450 2.4250 5.4350 2.4800 ;
	    RECT 0.5850 2.2500 5.4350 2.4250 ;
	    RECT 0.5850 2.1950 0.8750 2.2500 ;
	    RECT 2.3850 2.1950 2.6750 2.2500 ;
	    RECT 5.1450 2.1950 5.4350 2.2500 ;
	    RECT 5.1850 1.5750 5.4750 1.6300 ;
	    RECT 2.9200 1.4000 5.4750 1.5750 ;
	    RECT 2.9200 1.2050 3.1350 1.4000 ;
	    RECT 5.1850 1.3450 5.4750 1.4000 ;
	    RECT 1.0050 1.1500 1.2950 1.2050 ;
	    RECT 2.8450 1.1500 3.1350 1.2050 ;
	    RECT 1.0050 0.9750 3.1350 1.1500 ;
	    RECT 1.0050 0.9200 1.2950 0.9750 ;
	    RECT 2.8450 0.9200 3.1350 0.9750 ;
   END
END efs8hd_dfsbp_2
MACRO efs8hd_dfstp_2
   CLASS CORE ;
   FOREIGN efs8hd_dfstp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 9.6600 BY 3.4000 ;
   SITE unitehd ;
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 8.8100 2.0200 9.1400 3.0750 ;
	    RECT 8.8100 1.8700 9.5750 2.0200 ;
	    RECT 8.9750 1.8050 9.5750 1.8700 ;
	    RECT 9.0200 1.1200 9.5750 1.8050 ;
	    RECT 8.9900 1.0700 9.5750 1.1200 ;
	    RECT 8.9750 1.0300 9.5750 1.0700 ;
	    RECT 8.8900 0.9550 9.5750 1.0300 ;
	    RECT 8.8900 0.3300 9.1350 0.9550 ;
      END
   END Q
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.7700 1.2550 2.1800 2.0300 ;
      END
   END D
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 9.6600 3.5050 ;
	    RECT 0.5150 2.6700 0.8450 3.2950 ;
	    RECT 1.4550 2.6700 1.7850 3.2950 ;
	    RECT 3.4300 2.8200 3.8100 3.2950 ;
	    RECT 4.3300 2.8200 4.6600 3.2950 ;
	    RECT 5.9200 2.8200 6.3400 3.2950 ;
	    RECT 7.0100 2.4300 7.3400 3.2950 ;
	    RECT 8.4700 1.8700 8.6400 3.2950 ;
	    RECT 9.3100 2.2300 9.5750 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 9.6600 3.7000 ;
      END
   END vpwr
   PIN SETB
      PORT
         LAYER li1 ;
	    RECT 3.6100 0.9200 4.0200 1.3300 ;
	    RECT 6.6600 1.2550 7.0100 1.3300 ;
	    RECT 6.6600 0.9200 7.3400 1.2550 ;
         LAYER met1 ;
	    RECT 3.7650 1.1500 4.0550 1.2050 ;
	    RECT 6.9850 1.1500 7.2750 1.2050 ;
	    RECT 3.7650 0.9750 7.2750 1.1500 ;
	    RECT 3.7650 0.9200 4.0550 0.9750 ;
	    RECT 6.9850 0.9200 7.2750 0.9750 ;
      END
   END SETB
   PIN CLK
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.2200 0.4350 2.0300 ;
      END
   END CLK
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.4550 0.1050 1.7850 0.5800 ;
	    RECT 3.6100 0.1050 4.0200 0.6550 ;
	    RECT 4.7600 0.1050 5.0800 0.6800 ;
	    RECT 6.6900 0.1050 7.3300 0.7050 ;
	    RECT 8.3900 0.1050 8.7200 1.0300 ;
	    RECT 9.3050 0.1050 9.5750 0.7450 ;
	    RECT 0.0000 -0.1050 9.6600 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 9.6600 0.3000 ;
      END
   END vgnd
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.4550 0.3450 3.0800 ;
	    RECT 1.0150 2.5550 1.2350 3.0800 ;
	    RECT 0.0850 2.2450 0.8350 2.4550 ;
	    RECT 0.6050 1.0050 0.8350 2.2450 ;
	    RECT 0.0850 0.7950 0.8350 1.0050 ;
	    RECT 0.0850 0.4300 0.3450 0.7950 ;
	    RECT 1.0050 0.7050 1.2350 2.5550 ;
	    RECT 1.9550 2.4550 2.1250 3.0800 ;
	    RECT 2.3600 2.8150 3.1900 3.0250 ;
	    RECT 1.4300 2.2450 2.1250 2.4550 ;
	    RECT 1.4300 1.0300 1.6000 2.2450 ;
	    RECT 2.3500 1.9700 2.8500 2.4450 ;
	    RECT 1.4300 0.7950 2.1250 1.0300 ;
	    RECT 2.3500 0.8800 2.5700 1.9700 ;
	    RECT 3.0200 1.7550 3.1900 2.8150 ;
	    RECT 3.9900 2.6050 4.1600 2.9700 ;
	    RECT 5.1100 2.7050 5.7400 3.0200 ;
	    RECT 5.5700 2.6050 5.7400 2.7050 ;
	    RECT 6.5400 2.6050 6.7800 2.9700 ;
	    RECT 3.3600 2.2950 4.7100 2.6050 ;
	    RECT 3.3600 1.9700 3.6100 2.2950 ;
	    RECT 4.1200 1.7550 4.3700 1.9550 ;
	    RECT 3.0200 1.5450 4.3700 1.7550 ;
	    RECT 3.0200 1.4950 3.4400 1.5450 ;
	    RECT 2.7500 0.8050 3.1000 1.2700 ;
	    RECT 1.0150 0.4300 1.2350 0.7050 ;
	    RECT 1.9550 0.3800 2.1250 0.7950 ;
	    RECT 3.2700 0.5800 3.4400 1.4950 ;
	    RECT 4.5400 1.3300 4.7100 2.2950 ;
	    RECT 2.4250 0.3300 3.4400 0.5800 ;
	    RECT 4.3100 0.9050 4.7100 1.3300 ;
	    RECT 4.8800 2.0700 5.4000 2.4550 ;
	    RECT 5.5700 2.3950 6.7800 2.6050 ;
	    RECT 4.8800 1.1200 5.0500 2.0700 ;
	    RECT 5.2200 1.3300 5.4000 1.8450 ;
	    RECT 5.5700 1.7550 5.7400 2.3950 ;
	    RECT 7.5100 2.2050 7.6800 2.9700 ;
	    RECT 7.9700 2.3950 8.3000 3.0300 ;
	    RECT 7.5100 2.1800 7.8800 2.2050 ;
	    RECT 5.9100 1.9700 7.8800 2.1800 ;
	    RECT 5.5700 1.5450 7.4900 1.7550 ;
	    RECT 5.8000 1.1200 6.1500 1.2700 ;
	    RECT 4.8800 0.9050 6.1500 1.1200 ;
	    RECT 4.3100 0.3700 4.5600 0.9050 ;
	    RECT 6.3200 0.5950 6.4900 1.5450 ;
	    RECT 7.1400 1.4700 7.4900 1.5450 ;
	    RECT 7.6900 0.8500 7.8800 1.9700 ;
	    RECT 5.6400 0.3800 6.4900 0.5950 ;
	    RECT 7.5300 0.4400 7.8800 0.8500 ;
	    RECT 8.0500 1.6550 8.3000 2.3950 ;
	    RECT 8.0500 1.2450 8.8500 1.6550 ;
	    RECT 8.0500 0.4300 8.2200 1.2450 ;
         LAYER met1 ;
	    RECT 0.5450 2.4250 0.8350 2.4800 ;
	    RECT 2.3850 2.4250 2.6750 2.4800 ;
	    RECT 5.1450 2.4250 5.4350 2.4800 ;
	    RECT 0.5450 2.2500 5.4350 2.4250 ;
	    RECT 0.5450 2.1950 0.8350 2.2500 ;
	    RECT 2.3850 2.1950 2.6750 2.2500 ;
	    RECT 5.1450 2.1950 5.4350 2.2500 ;
	    RECT 5.1650 1.5750 5.4550 1.6300 ;
	    RECT 2.9200 1.4000 5.4550 1.5750 ;
	    RECT 2.9200 1.2050 3.1350 1.4000 ;
	    RECT 5.1650 1.3450 5.4550 1.4000 ;
	    RECT 1.0050 1.1500 1.2950 1.2050 ;
	    RECT 2.8450 1.1500 3.1350 1.2050 ;
	    RECT 1.0050 0.9750 3.1350 1.1500 ;
	    RECT 1.0050 0.9200 1.2950 0.9750 ;
	    RECT 2.8450 0.9200 3.1350 0.9750 ;
   END
END efs8hd_dfstp_2
MACRO efs8hd_dfxbp_2
   CLASS CORE ;
   FOREIGN efs8hd_dfxbp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 9.6600 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.4550 0.1050 1.7050 0.6800 ;
	    RECT 3.4000 0.1050 3.7700 0.7300 ;
	    RECT 5.5850 0.1050 5.7950 0.7700 ;
	    RECT 6.5600 0.1050 6.7300 0.8700 ;
	    RECT 7.4000 0.1050 7.5700 0.7500 ;
	    RECT 8.3900 0.1050 8.7200 1.0300 ;
	    RECT 9.3150 0.1050 9.5650 1.1300 ;
	    RECT 0.0000 -0.1050 9.6600 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 9.6600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 9.6600 3.5050 ;
	    RECT 0.5150 2.6700 0.8450 3.2950 ;
	    RECT 1.4400 2.7200 1.7050 3.2950 ;
	    RECT 3.6100 2.2950 3.7800 3.2950 ;
	    RECT 5.4900 2.6700 5.8050 3.2950 ;
	    RECT 6.5500 2.0300 6.7200 3.2950 ;
	    RECT 7.3900 2.1500 7.5650 3.2950 ;
	    RECT 8.4250 1.8700 8.6400 3.2950 ;
	    RECT 9.3150 1.8700 9.5650 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 9.6600 3.7000 ;
      END
   END vpwr
   PIN QN
      PORT
         LAYER li1 ;
	    RECT 8.8100 1.8700 9.1450 3.0800 ;
	    RECT 8.9300 1.1050 9.1450 1.8700 ;
	    RECT 8.8900 0.3300 9.1450 1.1050 ;
      END
   END QN
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.3700 0.8950 1.6500 2.0800 ;
      END
   END D
   PIN CLK
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.2200 0.4400 2.0300 ;
      END
   END CLK
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 6.8900 1.9700 7.2200 3.0250 ;
	    RECT 6.8900 1.8700 7.3000 1.9700 ;
	    RECT 7.0650 1.8050 7.3000 1.8700 ;
	    RECT 7.1100 1.0800 7.3000 1.8050 ;
	    RECT 7.0550 1.0300 7.3000 1.0800 ;
	    RECT 6.9000 0.9250 7.3000 1.0300 ;
	    RECT 6.9000 0.3800 7.2300 0.9250 ;
      END
   END Q
   OBS
         LAYER li1 ;
	    RECT 0.1750 2.4550 0.3450 3.0800 ;
	    RECT 0.1750 2.2450 0.8400 2.4550 ;
	    RECT 0.6100 1.0050 0.8400 2.2450 ;
	    RECT 0.1750 0.7950 0.8400 1.0050 ;
	    RECT 0.1750 0.4300 0.3450 0.7950 ;
	    RECT 1.0150 0.4300 1.2000 3.0800 ;
	    RECT 1.8750 2.5500 2.1250 3.0800 ;
	    RECT 2.3350 2.7400 3.4400 2.9500 ;
	    RECT 1.8200 2.3900 2.1250 2.5500 ;
	    RECT 1.8200 1.0050 1.9900 2.3900 ;
	    RECT 2.1600 1.4050 2.4000 2.1500 ;
	    RECT 2.5700 2.0700 3.1000 2.5250 ;
	    RECT 2.5700 1.1950 2.7400 2.0700 ;
	    RECT 3.2700 1.9700 3.4400 2.7400 ;
	    RECT 3.9500 2.6700 4.2000 3.0800 ;
	    RECT 4.4250 2.7050 5.3100 2.9200 ;
	    RECT 3.2700 1.8550 3.7800 1.9700 ;
	    RECT 1.8200 0.8450 2.0450 1.0050 ;
	    RECT 2.2150 0.9200 2.7400 1.1950 ;
	    RECT 2.9100 1.6450 3.7800 1.8550 ;
	    RECT 1.8750 0.6700 2.0450 0.8450 ;
	    RECT 2.9100 0.6700 3.0800 1.6450 ;
	    RECT 3.6100 1.5550 3.7800 1.6450 ;
	    RECT 3.2900 1.3300 3.4900 1.3700 ;
	    RECT 3.9500 1.3300 4.1200 2.6700 ;
	    RECT 4.2900 1.5550 4.4800 2.4550 ;
	    RECT 3.2900 0.9550 4.1200 1.3300 ;
	    RECT 4.6500 1.2950 4.9700 2.4950 ;
	    RECT 1.8750 0.4550 2.2100 0.6700 ;
	    RECT 2.4050 0.4550 3.0800 0.6700 ;
	    RECT 3.9500 0.6700 4.1200 0.9550 ;
	    RECT 4.5050 0.8800 4.9700 1.2950 ;
	    RECT 5.1400 1.6550 5.3100 2.7050 ;
	    RECT 6.0400 2.3800 6.3800 3.0800 ;
	    RECT 5.4800 1.9150 6.3800 2.3800 ;
	    RECT 7.9050 2.1450 8.2350 3.0550 ;
	    RECT 6.1900 1.6550 6.3800 1.9150 ;
	    RECT 7.9650 1.6550 8.2350 2.1450 ;
	    RECT 5.1400 1.2450 6.0200 1.6550 ;
	    RECT 6.1900 1.2450 6.9400 1.6550 ;
	    RECT 7.9650 1.2450 8.7600 1.6550 ;
	    RECT 5.1400 0.6700 5.3100 1.2450 ;
	    RECT 6.1900 1.0300 6.3900 1.2450 ;
	    RECT 3.9500 0.4550 4.3550 0.6700 ;
	    RECT 4.5250 0.4550 5.3100 0.6700 ;
	    RECT 6.0600 0.3750 6.3900 1.0300 ;
	    RECT 7.9650 0.7700 8.1650 1.2450 ;
	    RECT 7.9050 0.4300 8.1650 0.7700 ;
         LAYER met1 ;
	    RECT 0.5700 2.4250 0.8600 2.4800 ;
	    RECT 2.6700 2.4250 2.9600 2.4800 ;
	    RECT 4.2400 2.4250 4.5300 2.4800 ;
	    RECT 0.5700 2.2500 4.5300 2.4250 ;
	    RECT 0.5700 2.1950 0.8600 2.2500 ;
	    RECT 2.6700 2.1950 2.9600 2.2500 ;
	    RECT 4.2400 2.1950 4.5300 2.2500 ;
	    RECT 0.9650 2.0000 1.2550 2.0550 ;
	    RECT 2.1550 2.0000 2.4450 2.0550 ;
	    RECT 4.6750 2.0000 4.9650 2.0550 ;
	    RECT 0.9650 1.8250 4.9650 2.0000 ;
	    RECT 0.9650 1.7700 1.2550 1.8250 ;
	    RECT 2.1550 1.7700 2.4450 1.8250 ;
	    RECT 4.6750 1.7700 4.9650 1.8250 ;
   END
END efs8hd_dfxbp_2
MACRO efs8hd_dfxtp_2
   CLASS CORE ;
   FOREIGN efs8hd_dfxtp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 7.8200 BY 3.4000 ;
   SITE unitehd ;
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 6.8850 1.9700 7.2150 3.0250 ;
	    RECT 6.8850 1.8700 7.2750 1.9700 ;
	    RECT 7.0600 1.8050 7.2750 1.8700 ;
	    RECT 7.1050 1.0800 7.2750 1.8050 ;
	    RECT 7.0500 1.0300 7.2750 1.0800 ;
	    RECT 6.8950 0.9250 7.2750 1.0300 ;
	    RECT 6.8950 0.3800 7.2250 0.9250 ;
      END
   END Q
   PIN CLK
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.2200 0.4400 2.0300 ;
      END
   END CLK
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.3700 0.8950 1.6500 2.0800 ;
      END
   END D
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 7.8200 3.5050 ;
	    RECT 0.5150 2.6700 0.8450 3.2950 ;
	    RECT 1.4400 2.7200 1.7050 3.2950 ;
	    RECT 3.6100 2.2950 3.7800 3.2950 ;
	    RECT 5.4900 2.6700 5.8050 3.2950 ;
	    RECT 6.5450 2.0300 6.7150 3.2950 ;
	    RECT 7.3850 2.1500 7.5550 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 7.8200 3.7000 ;
      END
   END vpwr
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.4550 0.1050 1.7050 0.6800 ;
	    RECT 3.4000 0.1050 3.7700 0.7300 ;
	    RECT 5.5850 0.1050 5.7950 0.7700 ;
	    RECT 6.5550 0.1050 6.7250 0.8700 ;
	    RECT 7.3950 0.1050 7.5650 0.7500 ;
	    RECT 0.0000 -0.1050 7.8200 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 7.8200 0.3000 ;
      END
   END vgnd
   OBS
         LAYER li1 ;
	    RECT 0.1750 2.4550 0.3450 3.0800 ;
	    RECT 0.1750 2.2450 0.8400 2.4550 ;
	    RECT 0.6100 1.0050 0.8400 2.2450 ;
	    RECT 0.1750 0.7950 0.8400 1.0050 ;
	    RECT 0.1750 0.4300 0.3450 0.7950 ;
	    RECT 1.0150 0.4300 1.2000 3.0800 ;
	    RECT 1.8750 2.5500 2.1250 3.0800 ;
	    RECT 2.3350 2.7400 3.4400 2.9500 ;
	    RECT 1.8200 2.3900 2.1250 2.5500 ;
	    RECT 1.8200 1.0050 1.9900 2.3900 ;
	    RECT 2.1600 1.4050 2.4000 2.1500 ;
	    RECT 2.5700 2.0700 3.1000 2.5250 ;
	    RECT 2.5700 1.1950 2.7400 2.0700 ;
	    RECT 3.2700 1.9700 3.4400 2.7400 ;
	    RECT 3.9500 2.6700 4.2000 3.0800 ;
	    RECT 4.4250 2.7050 5.3100 2.9200 ;
	    RECT 3.2700 1.8550 3.7800 1.9700 ;
	    RECT 1.8200 0.8450 2.0450 1.0050 ;
	    RECT 2.2150 0.9200 2.7400 1.1950 ;
	    RECT 2.9100 1.6450 3.7800 1.8550 ;
	    RECT 1.8750 0.6700 2.0450 0.8450 ;
	    RECT 2.9100 0.6700 3.0800 1.6450 ;
	    RECT 3.6100 1.5550 3.7800 1.6450 ;
	    RECT 3.2900 1.3300 3.4900 1.3700 ;
	    RECT 3.9500 1.3300 4.1200 2.6700 ;
	    RECT 4.2900 1.5550 4.4800 2.4550 ;
	    RECT 3.2900 0.9550 4.1200 1.3300 ;
	    RECT 4.6500 1.2950 4.9700 2.4950 ;
	    RECT 1.8750 0.4550 2.2100 0.6700 ;
	    RECT 2.4050 0.4550 3.0800 0.6700 ;
	    RECT 3.9500 0.6700 4.1200 0.9550 ;
	    RECT 4.5050 0.8800 4.9700 1.2950 ;
	    RECT 5.1400 1.6550 5.3100 2.7050 ;
	    RECT 6.0350 2.3800 6.3750 3.0800 ;
	    RECT 5.4800 1.9150 6.3750 2.3800 ;
	    RECT 6.1850 1.6550 6.3750 1.9150 ;
	    RECT 5.1400 1.2450 6.0150 1.6550 ;
	    RECT 6.1850 1.2450 6.9350 1.6550 ;
	    RECT 5.1400 0.6700 5.3100 1.2450 ;
	    RECT 6.1850 1.0300 6.3850 1.2450 ;
	    RECT 3.9500 0.4550 4.3550 0.6700 ;
	    RECT 4.5250 0.4550 5.3100 0.6700 ;
	    RECT 6.0550 0.3750 6.3850 1.0300 ;
         LAYER met1 ;
	    RECT 0.5700 2.4250 0.8600 2.4800 ;
	    RECT 2.6700 2.4250 2.9600 2.4800 ;
	    RECT 4.2400 2.4250 4.5300 2.4800 ;
	    RECT 0.5700 2.2500 4.5300 2.4250 ;
	    RECT 0.5700 2.1950 0.8600 2.2500 ;
	    RECT 2.6700 2.1950 2.9600 2.2500 ;
	    RECT 4.2400 2.1950 4.5300 2.2500 ;
	    RECT 0.9650 2.0000 1.2550 2.0550 ;
	    RECT 2.1550 2.0000 2.4450 2.0550 ;
	    RECT 4.6750 2.0000 4.9650 2.0550 ;
	    RECT 0.9650 1.8250 4.9650 2.0000 ;
	    RECT 0.9650 1.7700 1.2550 1.8250 ;
	    RECT 2.1550 1.7700 2.4450 1.8250 ;
	    RECT 4.6750 1.7700 4.9650 1.8250 ;
   END
END efs8hd_dfxtp_2
MACRO efs8hd_dlclkp_2
   CLASS CORE ;
   FOREIGN efs8hd_dlclkp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 6.9000 BY 3.4000 ;
   SITE unitehd ;
   PIN GATE
      PORT
         LAYER li1 ;
	    RECT 1.5300 1.7950 2.2150 2.1050 ;
	    RECT 1.9850 0.3550 2.2150 1.7950 ;
      END
   END GATE
   PIN GCLK
      PORT
         LAYER li1 ;
	    RECT 6.0950 1.8700 6.3600 3.0700 ;
	    RECT 6.1650 0.7450 6.3600 1.8700 ;
	    RECT 6.0600 0.3200 6.3600 0.7450 ;
      END
   END GCLK
   PIN CLK
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.2300 0.3300 2.0300 ;
	    RECT 5.2100 1.3800 5.4850 1.7950 ;
         LAYER met1 ;
	    RECT 0.0900 1.5750 0.3800 1.6300 ;
	    RECT 5.1500 1.5750 5.4400 1.6300 ;
	    RECT 0.0900 1.4000 5.4400 1.5750 ;
	    RECT 0.0900 1.3450 0.3800 1.4000 ;
	    RECT 5.1500 1.3450 5.4400 1.4000 ;
      END
   END CLK
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5550 ;
	    RECT 1.4850 0.1050 1.8150 1.1300 ;
	    RECT 3.8950 0.1050 4.1450 0.7650 ;
	    RECT 5.6750 0.1050 5.8450 0.6800 ;
	    RECT 6.5300 0.1050 6.8100 1.1050 ;
	    RECT 0.0000 -0.1050 6.9000 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 6.9000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 6.9000 3.5050 ;
	    RECT 0.5150 2.6700 0.8450 3.2950 ;
	    RECT 1.4550 2.7450 1.8200 3.2950 ;
	    RECT 3.4000 2.6700 3.7000 3.2950 ;
	    RECT 4.3150 2.5150 4.6000 3.2950 ;
	    RECT 5.5750 2.6650 5.9250 3.2950 ;
	    RECT 6.5300 1.8550 6.8100 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 6.9000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1750 2.4550 0.3450 3.0800 ;
	    RECT 1.0150 2.5300 1.2400 3.0800 ;
	    RECT 2.4800 2.8200 3.2300 3.0300 ;
	    RECT 0.1750 2.2450 0.7800 2.4550 ;
	    RECT 0.6100 1.7400 0.7800 2.2450 ;
	    RECT 1.0150 2.3200 2.6450 2.5300 ;
	    RECT 0.6100 1.3250 0.8400 1.7400 ;
	    RECT 0.6100 0.9800 0.7800 1.3250 ;
	    RECT 0.1750 0.7700 0.7800 0.9800 ;
	    RECT 0.1750 0.3250 0.3450 0.7700 ;
	    RECT 1.0150 0.3250 1.2800 2.3200 ;
	    RECT 2.3950 1.2300 2.6450 2.3200 ;
	    RECT 3.0600 1.6550 3.2300 2.8200 ;
	    RECT 3.9150 2.3300 4.1350 3.0450 ;
	    RECT 3.4350 2.3000 4.1350 2.3300 ;
	    RECT 5.0100 2.3700 5.3400 3.0800 ;
	    RECT 3.4350 1.9200 4.7350 2.3000 ;
	    RECT 5.0100 2.1550 5.9250 2.3700 ;
	    RECT 3.0600 1.4450 4.1800 1.6550 ;
	    RECT 3.5550 1.2450 4.1800 1.4450 ;
	    RECT 4.3500 1.2450 4.7350 1.9200 ;
	    RECT 5.7550 1.6550 5.9250 2.1550 ;
	    RECT 2.3950 1.0200 3.2250 1.2300 ;
	    RECT 3.5550 0.7000 3.7250 1.2450 ;
	    RECT 4.3500 0.7700 4.5850 1.2450 ;
	    RECT 5.7550 1.1700 5.9950 1.6550 ;
	    RECT 4.9300 0.9550 5.9950 1.1700 ;
	    RECT 4.9300 0.7750 5.1500 0.9550 ;
	    RECT 2.7950 0.4900 3.7250 0.7000 ;
	    RECT 4.3150 0.3200 4.5850 0.7700 ;
	    RECT 4.8350 0.3650 5.1500 0.7750 ;
   END
END efs8hd_dlclkp_2
MACRO efs8hd_dlrbp_2
   CLASS CORE ;
   FOREIGN efs8hd_dlrbp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 8.2800 BY 3.4000 ;
   SITE unitehd ;
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 5.6800 2.0750 5.9300 3.0800 ;
	    RECT 5.6800 1.8700 6.0650 2.0750 ;
	    RECT 5.7900 1.6550 6.0650 1.8700 ;
	    RECT 5.7900 1.1050 6.3600 1.6550 ;
	    RECT 5.7900 1.0450 6.1500 1.1050 ;
	    RECT 5.6800 0.8300 6.1500 1.0450 ;
	    RECT 5.6800 0.4150 5.8500 0.8300 ;
      END
   END Q
   PIN RESETB
      PORT
         LAYER li1 ;
	    RECT 4.4000 1.2450 5.1500 1.6550 ;
      END
   END RESETB
   PIN QN
      PORT
         LAYER li1 ;
	    RECT 7.5150 2.0050 7.7650 3.0800 ;
	    RECT 7.5950 1.6550 7.7650 2.0050 ;
	    RECT 7.5950 1.3200 8.1950 1.6550 ;
	    RECT 7.5950 1.0300 7.7650 1.3200 ;
	    RECT 7.5150 0.3200 7.7650 1.0300 ;
      END
   END QN
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.4600 1.1950 1.7900 1.6550 ;
      END
   END D
   PIN GATE
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.2300 0.3300 2.0300 ;
      END
   END GATE
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.8750 0.1050 2.2050 0.5550 ;
	    RECT 3.7400 0.1050 4.0700 0.6650 ;
	    RECT 5.1100 0.1050 5.4900 0.6050 ;
	    RECT 6.0200 0.1050 6.3600 0.5800 ;
	    RECT 7.0350 0.1050 7.3400 0.6800 ;
	    RECT 7.9350 0.1050 8.1950 1.1050 ;
	    RECT 0.0000 -0.1050 8.2800 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 8.2800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 8.2800 3.5050 ;
	    RECT 0.5150 2.6700 0.8450 3.2950 ;
	    RECT 1.9550 2.2950 2.2700 3.2950 ;
	    RECT 3.7550 2.6700 4.6000 3.2950 ;
	    RECT 5.1100 2.3450 5.4900 3.2950 ;
	    RECT 6.1000 2.2900 6.3600 3.2950 ;
	    RECT 7.0450 2.2950 7.3400 3.2950 ;
	    RECT 7.9350 1.8700 8.1950 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 8.2800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.4550 0.3450 3.0800 ;
	    RECT 0.0850 2.2450 0.7800 2.4550 ;
	    RECT 0.6100 1.7500 0.7800 2.2450 ;
	    RECT 1.0150 2.1050 1.2400 3.0800 ;
	    RECT 0.6100 1.3400 0.8400 1.7500 ;
	    RECT 0.6100 1.0050 0.7800 1.3400 ;
	    RECT 0.0850 0.7950 0.7800 1.0050 ;
	    RECT 0.0850 0.4300 0.3450 0.7950 ;
	    RECT 1.0150 0.4300 1.1850 2.1050 ;
	    RECT 1.4550 2.0800 1.7850 3.0200 ;
	    RECT 2.7450 2.8200 3.5850 3.0300 ;
	    RECT 3.2700 2.6550 3.5850 2.8200 ;
	    RECT 3.3050 2.5950 3.5850 2.6550 ;
	    RECT 3.3950 2.5550 3.5850 2.5950 ;
	    RECT 3.3950 2.5200 3.6050 2.5550 ;
	    RECT 2.9250 2.3800 3.1250 2.4950 ;
	    RECT 3.4150 2.4900 3.6050 2.5200 ;
	    RECT 3.4200 2.4700 3.6050 2.4900 ;
	    RECT 3.4300 2.4500 3.6050 2.4700 ;
	    RECT 1.4550 1.8700 2.1400 2.0800 ;
	    RECT 1.9700 1.3700 2.1400 1.8700 ;
	    RECT 2.4700 1.6950 2.7550 2.1050 ;
	    RECT 2.9250 1.9700 3.2650 2.3800 ;
	    RECT 1.9700 0.9800 2.3400 1.3700 ;
	    RECT 2.9250 1.2950 3.0950 1.9700 ;
	    RECT 3.4350 1.6550 3.6050 2.4500 ;
	    RECT 4.7700 2.3300 4.9400 3.0450 ;
	    RECT 3.8400 2.1300 4.9400 2.3300 ;
	    RECT 3.8400 1.9200 5.5100 2.1300 ;
	    RECT 5.3200 1.6550 5.5100 1.9200 ;
	    RECT 6.5350 1.6550 6.8700 3.0800 ;
	    RECT 3.4350 1.4550 4.2000 1.6550 ;
	    RECT 1.5350 0.9550 2.3400 0.9800 ;
	    RECT 1.5350 0.7700 2.1400 0.9550 ;
	    RECT 2.7150 0.8800 3.0950 1.2950 ;
	    RECT 3.3300 1.2450 4.2000 1.4550 ;
	    RECT 5.3200 1.2450 5.6200 1.6550 ;
	    RECT 6.5350 1.2450 7.4250 1.6550 ;
	    RECT 1.5350 0.4300 1.7050 0.7700 ;
	    RECT 3.3300 0.6700 3.5000 1.2450 ;
	    RECT 5.3200 1.0300 5.5100 1.2450 ;
	    RECT 2.7700 0.4550 3.5000 0.6700 ;
	    RECT 4.2700 0.8200 5.5100 1.0300 ;
	    RECT 4.2700 0.5200 4.5700 0.8200 ;
	    RECT 6.5350 0.3200 6.8650 1.2450 ;
         LAYER met1 ;
	    RECT 1.0100 2.4250 1.3000 2.4800 ;
	    RECT 2.8700 2.4250 3.1600 2.4800 ;
	    RECT 1.0100 2.2500 3.1600 2.4250 ;
	    RECT 1.0100 2.1950 1.3000 2.2500 ;
	    RECT 2.8700 2.1950 3.1600 2.2500 ;
	    RECT 0.5500 2.0000 0.8400 2.0550 ;
	    RECT 2.4100 2.0000 2.7000 2.0550 ;
	    RECT 0.5500 1.8250 2.7000 2.0000 ;
	    RECT 0.5500 1.7700 0.8400 1.8250 ;
	    RECT 2.4100 1.7700 2.7000 1.8250 ;
   END
END efs8hd_dlrbp_2
MACRO efs8hd_dlrtn_2
   CLASS CORE ;
   FOREIGN efs8hd_dlrtn_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 6.4400 BY 3.4000 ;
   SITE unitehd ;
   PIN RESETB
      PORT
         LAYER li1 ;
	    RECT 4.4800 1.2450 5.1700 1.6550 ;
      END
   END RESETB
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 5.6550 2.3450 5.9250 3.0800 ;
	    RECT 5.7550 1.8750 5.9250 2.3450 ;
	    RECT 5.7550 1.7800 6.3550 1.8750 ;
	    RECT 5.7600 1.7700 6.3550 1.7800 ;
	    RECT 5.7650 1.7650 6.3550 1.7700 ;
	    RECT 5.7750 1.7300 6.3550 1.7650 ;
	    RECT 5.7850 1.1150 6.3550 1.7300 ;
	    RECT 5.7700 1.0800 6.3550 1.1150 ;
	    RECT 5.7550 0.9550 6.3550 1.0800 ;
	    RECT 5.7550 0.6050 5.9250 0.9550 ;
	    RECT 5.5950 0.3200 5.9250 0.6050 ;
      END
   END Q
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.4600 1.1950 1.7900 1.6550 ;
      END
   END D
   PIN GATEN
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.2300 0.3300 2.0300 ;
      END
   END GATEN
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.8750 0.1050 2.2050 0.5550 ;
	    RECT 3.7350 0.1050 4.0700 0.6650 ;
	    RECT 5.0950 0.1050 5.4250 0.6050 ;
	    RECT 6.0950 0.1050 6.3550 0.7450 ;
	    RECT 0.0000 -0.1050 6.4400 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 6.4400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 6.4400 3.5050 ;
	    RECT 0.5150 2.6700 0.8450 3.2950 ;
	    RECT 1.9550 2.2950 2.2700 3.2950 ;
	    RECT 3.8000 2.6700 4.1100 3.2950 ;
	    RECT 4.2800 2.6700 4.5600 3.2950 ;
	    RECT 5.0900 2.3450 5.4600 3.2950 ;
	    RECT 6.0950 2.0900 6.3550 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 6.4400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1750 2.4550 0.3450 3.0800 ;
	    RECT 0.1750 2.2450 0.7800 2.4550 ;
	    RECT 0.6100 1.7500 0.7800 2.2450 ;
	    RECT 1.0150 2.1050 1.2400 3.0800 ;
	    RECT 0.6100 1.3400 0.8400 1.7500 ;
	    RECT 0.6100 1.0050 0.7800 1.3400 ;
	    RECT 0.1750 0.7950 0.7800 1.0050 ;
	    RECT 0.1750 0.4300 0.3450 0.7950 ;
	    RECT 1.0150 0.4300 1.1850 2.1050 ;
	    RECT 1.4550 2.0800 1.7850 3.0200 ;
	    RECT 2.7750 2.8200 3.6050 3.0300 ;
	    RECT 1.4550 1.8700 2.1400 2.0800 ;
	    RECT 1.9600 1.3700 2.1400 1.8700 ;
	    RECT 2.4700 1.6950 2.7550 2.5050 ;
	    RECT 2.9250 1.7700 3.2650 2.4950 ;
	    RECT 2.9250 1.4300 3.0950 1.7700 ;
	    RECT 3.4350 1.6550 3.6050 2.8200 ;
	    RECT 4.7300 2.3300 4.9200 3.0800 ;
	    RECT 3.8200 2.1300 4.9200 2.3300 ;
	    RECT 3.8200 1.9200 5.5850 2.1300 ;
	    RECT 5.4150 1.6550 5.5850 1.9200 ;
	    RECT 3.4350 1.5550 4.3100 1.6550 ;
	    RECT 1.9600 0.9800 2.3400 1.3700 ;
	    RECT 1.5350 0.9550 2.3400 0.9800 ;
	    RECT 1.5350 0.7700 2.1400 0.9550 ;
	    RECT 2.6750 0.8800 3.0950 1.4300 ;
	    RECT 3.3300 1.2800 4.3100 1.5550 ;
	    RECT 1.5350 0.4300 1.7050 0.7700 ;
	    RECT 3.3300 0.6700 3.5000 1.2800 ;
	    RECT 5.3500 1.2450 5.6150 1.6550 ;
	    RECT 5.4150 1.0300 5.5850 1.2450 ;
	    RECT 2.8100 0.4550 3.5000 0.6700 ;
	    RECT 4.2400 0.8200 5.5850 1.0300 ;
	    RECT 4.2400 0.3200 4.5900 0.8200 ;
         LAYER met1 ;
	    RECT 1.0100 2.4250 1.3000 2.4800 ;
	    RECT 2.4100 2.4250 2.7000 2.4800 ;
	    RECT 1.0100 2.2500 2.7000 2.4250 ;
	    RECT 1.0100 2.1950 1.3000 2.2500 ;
	    RECT 2.4100 2.1950 2.7000 2.2500 ;
	    RECT 0.5500 2.0000 0.8400 2.0550 ;
	    RECT 2.8700 2.0000 3.1600 2.0550 ;
	    RECT 0.5500 1.8250 3.1600 2.0000 ;
	    RECT 0.5500 1.7700 0.8400 1.8250 ;
	    RECT 2.8700 1.7700 3.1600 1.8250 ;
   END
END efs8hd_dlrtn_2
MACRO efs8hd_dlrtp_2
   CLASS CORE ;
   FOREIGN efs8hd_dlrtp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 6.4400 BY 3.4000 ;
   SITE unitehd ;
   PIN RESETB
      PORT
         LAYER li1 ;
	    RECT 4.4800 1.2950 5.2400 1.6550 ;
	    RECT 4.4800 1.2450 4.8150 1.2950 ;
      END
   END RESETB
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 5.6550 2.3450 5.9250 3.0800 ;
	    RECT 5.7550 1.8750 5.9250 2.3450 ;
	    RECT 5.7550 1.7800 6.3550 1.8750 ;
	    RECT 5.7600 1.7700 6.3550 1.7800 ;
	    RECT 5.7650 1.7650 6.3550 1.7700 ;
	    RECT 5.7750 1.7300 6.3550 1.7650 ;
	    RECT 5.7850 1.1150 6.3550 1.7300 ;
	    RECT 5.7700 1.0800 6.3550 1.1150 ;
	    RECT 5.7550 0.9550 6.3550 1.0800 ;
	    RECT 5.7550 0.6050 5.9250 0.9550 ;
	    RECT 5.5950 0.3200 5.9250 0.6050 ;
      END
   END Q
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.4400 1.1950 1.7700 1.6550 ;
      END
   END D
   PIN GATE
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.2300 0.3300 2.0300 ;
      END
   END GATE
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.8750 0.1050 2.2050 0.5550 ;
	    RECT 3.7200 0.1050 4.0600 0.6650 ;
	    RECT 5.2550 0.1050 5.4250 0.6550 ;
	    RECT 6.0950 0.1050 6.3550 0.7450 ;
	    RECT 0.0000 -0.1050 6.4400 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 6.4400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 6.4400 3.5050 ;
	    RECT 0.5150 2.6700 0.8450 3.2950 ;
	    RECT 1.9550 2.2950 2.2500 3.2950 ;
	    RECT 3.7500 2.7200 4.0900 3.2950 ;
	    RECT 4.2800 2.6700 4.5600 3.2950 ;
	    RECT 5.1400 2.3450 5.4850 3.2950 ;
	    RECT 6.0950 2.0900 6.3550 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 6.4400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1750 2.4550 0.3450 3.0800 ;
	    RECT 0.1750 2.2450 0.7800 2.4550 ;
	    RECT 0.6100 1.7500 0.7800 2.2450 ;
	    RECT 1.0150 2.1050 1.2400 3.0800 ;
	    RECT 0.6100 1.3400 0.8400 1.7500 ;
	    RECT 0.6100 1.0050 0.7800 1.3400 ;
	    RECT 0.0850 0.7950 0.7800 1.0050 ;
	    RECT 0.0850 0.4300 0.3450 0.7950 ;
	    RECT 1.0150 0.4300 1.1850 2.1050 ;
	    RECT 1.4350 2.0800 1.7850 3.0200 ;
	    RECT 2.7700 2.8200 3.5800 3.0300 ;
	    RECT 3.4100 2.6050 3.5800 2.8200 ;
	    RECT 3.4100 2.5000 3.6050 2.6050 ;
	    RECT 3.4150 2.4950 3.6050 2.5000 ;
	    RECT 2.9050 2.3900 3.1750 2.4950 ;
	    RECT 3.4200 2.4800 3.6050 2.4950 ;
	    RECT 2.9050 2.2250 3.2650 2.3900 ;
	    RECT 1.4350 1.8700 2.1200 2.0800 ;
	    RECT 1.9500 1.3700 2.1200 1.8700 ;
	    RECT 2.4500 1.6950 2.7550 2.1050 ;
	    RECT 2.9300 1.9650 3.2650 2.2250 ;
	    RECT 1.9500 0.9800 2.3350 1.3700 ;
	    RECT 2.9300 1.3000 3.1000 1.9650 ;
	    RECT 3.4350 1.6550 3.6050 2.4800 ;
	    RECT 4.8000 2.3300 4.9700 3.0800 ;
	    RECT 3.7750 2.1300 4.9700 2.3300 ;
	    RECT 3.7750 1.9200 5.5850 2.1300 ;
	    RECT 5.4150 1.6550 5.5850 1.9200 ;
	    RECT 1.5150 0.9550 2.3350 0.9800 ;
	    RECT 1.5150 0.7700 2.1200 0.9550 ;
	    RECT 2.5850 0.9200 3.1000 1.3000 ;
	    RECT 3.2700 1.2450 4.2200 1.6550 ;
	    RECT 5.4150 1.2450 5.6150 1.6550 ;
	    RECT 1.5150 0.4300 1.7050 0.7700 ;
	    RECT 3.2700 0.6700 3.4450 1.2450 ;
	    RECT 5.4150 1.0800 5.5850 1.2450 ;
	    RECT 4.9550 1.0300 5.5850 1.0800 ;
	    RECT 2.7700 0.4550 3.4450 0.6700 ;
	    RECT 4.2400 0.8700 5.5850 1.0300 ;
	    RECT 4.2400 0.8200 5.0950 0.8700 ;
	    RECT 4.2400 0.3200 4.5800 0.8200 ;
         LAYER met1 ;
	    RECT 1.0100 2.4250 1.3000 2.4800 ;
	    RECT 2.8650 2.4250 3.1550 2.4800 ;
	    RECT 1.0100 2.2500 3.1550 2.4250 ;
	    RECT 1.0100 2.1950 1.3000 2.2500 ;
	    RECT 2.8650 2.1950 3.1550 2.2500 ;
	    RECT 0.5500 2.0000 0.8400 2.0550 ;
	    RECT 2.3900 2.0000 2.6800 2.0550 ;
	    RECT 0.5500 1.8250 2.6800 2.0000 ;
	    RECT 0.5500 1.7700 0.8400 1.8250 ;
	    RECT 2.3900 1.7700 2.6800 1.8250 ;
   END
END efs8hd_dlrtp_2
MACRO efs8hd_dlxbn_2
   CLASS CORE ;
   FOREIGN efs8hd_dlxbn_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 7.8200 BY 3.4000 ;
   SITE unitehd ;
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.4800 1.1950 1.8100 1.6550 ;
      END
   END D
   PIN GATEN
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.2300 0.3300 2.0300 ;
      END
   END GATEN
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 5.2150 2.1400 5.4650 3.0700 ;
	    RECT 5.2150 1.8700 5.5000 2.1400 ;
	    RECT 5.3300 1.6550 5.5000 1.8700 ;
	    RECT 5.3300 1.2450 5.9050 1.6550 ;
	    RECT 5.3300 1.0300 5.5000 1.2450 ;
	    RECT 5.2150 0.8250 5.5000 1.0300 ;
	    RECT 5.2150 0.5200 5.4650 0.8250 ;
      END
   END Q
   PIN QN
      PORT
         LAYER li1 ;
	    RECT 7.0500 1.8050 7.3050 3.0800 ;
	    RECT 7.0950 1.6550 7.3050 1.8050 ;
	    RECT 7.0950 1.3200 7.7350 1.6550 ;
	    RECT 7.0950 1.0300 7.3050 1.3200 ;
	    RECT 7.0500 0.3200 7.3050 1.0300 ;
      END
   END QN
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 7.8200 3.5050 ;
	    RECT 0.5150 2.6700 0.8450 3.2950 ;
	    RECT 1.9750 2.2950 2.2900 3.2950 ;
	    RECT 3.8400 2.6700 4.1400 3.2950 ;
	    RECT 4.7600 1.8700 5.0450 3.2950 ;
	    RECT 5.6350 2.2950 5.9050 3.2950 ;
	    RECT 6.5850 2.2950 6.8800 3.2950 ;
	    RECT 7.4750 1.8700 7.7350 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 7.8200 3.7000 ;
      END
   END vpwr
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.8950 0.1050 2.2250 0.5550 ;
	    RECT 3.7600 0.1050 4.0900 1.0300 ;
	    RECT 4.7600 0.1050 5.0450 1.0300 ;
	    RECT 5.6350 0.1050 5.9050 0.6800 ;
	    RECT 6.5850 0.1050 6.8800 0.6800 ;
	    RECT 7.4750 0.1050 7.7350 1.1050 ;
	    RECT 0.0000 -0.1050 7.8200 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 7.8200 0.3000 ;
      END
   END vgnd
   OBS
         LAYER li1 ;
	    RECT 0.1750 2.4550 0.3450 3.0800 ;
	    RECT 0.1750 2.2450 0.7800 2.4550 ;
	    RECT 0.6100 1.7500 0.7800 2.2450 ;
	    RECT 1.0150 2.1050 1.2400 3.0800 ;
	    RECT 0.6100 1.3400 0.8400 1.7500 ;
	    RECT 0.6100 1.0050 0.7800 1.3400 ;
	    RECT 0.1750 0.7950 0.7800 1.0050 ;
	    RECT 0.1750 0.4300 0.3450 0.7950 ;
	    RECT 1.0150 0.4300 1.1850 2.1050 ;
	    RECT 1.4750 2.0800 1.8050 3.0200 ;
	    RECT 2.9200 2.8200 3.6700 3.0300 ;
	    RECT 1.4750 1.8700 2.1600 2.0800 ;
	    RECT 1.9900 1.3700 2.1600 1.8700 ;
	    RECT 2.4900 1.6950 2.7750 2.5050 ;
	    RECT 2.9450 1.7700 3.2850 2.4950 ;
	    RECT 1.9900 0.9800 2.3600 1.3700 ;
	    RECT 2.9450 1.2950 3.1150 1.7700 ;
	    RECT 3.5000 1.6550 3.6700 2.8200 ;
	    RECT 4.3600 2.3300 4.5800 3.0450 ;
	    RECT 3.8600 1.9200 4.5800 2.3300 ;
	    RECT 4.4100 1.6550 4.5800 1.9200 ;
	    RECT 6.0750 1.6550 6.4050 3.0800 ;
	    RECT 3.5000 1.4550 4.2200 1.6550 ;
	    RECT 1.5550 0.9550 2.3600 0.9800 ;
	    RECT 1.5550 0.7700 2.1600 0.9550 ;
	    RECT 2.7350 0.8800 3.1150 1.2950 ;
	    RECT 3.3500 1.2450 4.2200 1.4550 ;
	    RECT 4.4100 1.2450 5.1600 1.6550 ;
	    RECT 6.0750 1.2450 6.9250 1.6550 ;
	    RECT 1.5550 0.4300 1.7250 0.7700 ;
	    RECT 3.3500 0.6700 3.5200 1.2450 ;
	    RECT 4.4100 1.0300 4.5800 1.2450 ;
	    RECT 2.8600 0.4550 3.5200 0.6700 ;
	    RECT 4.3600 0.5200 4.5800 1.0300 ;
	    RECT 6.0750 0.3200 6.4050 1.2450 ;
         LAYER met1 ;
	    RECT 1.0100 2.4250 1.3000 2.4800 ;
	    RECT 2.4300 2.4250 2.7200 2.4800 ;
	    RECT 1.0100 2.2500 2.7200 2.4250 ;
	    RECT 1.0100 2.1950 1.3000 2.2500 ;
	    RECT 2.4300 2.1950 2.7200 2.2500 ;
	    RECT 0.5500 2.0000 0.8400 2.0550 ;
	    RECT 2.8900 2.0000 3.1800 2.0550 ;
	    RECT 0.5500 1.8250 3.1800 2.0000 ;
	    RECT 0.5500 1.7700 0.8400 1.8250 ;
	    RECT 2.8900 1.7700 3.1800 1.8250 ;
   END
END efs8hd_dlxbn_2
MACRO efs8hd_dlxtn_2
   CLASS CORE ;
   FOREIGN efs8hd_dlxtn_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.9800 BY 3.4000 ;
   SITE unitehd ;
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.4800 1.1950 1.8100 1.6550 ;
      END
   END D
   PIN GATEN
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.2300 0.3300 2.0300 ;
      END
   END GATEN
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 5.2150 2.0500 5.4650 3.0700 ;
	    RECT 5.2150 1.8700 5.5000 2.0500 ;
	    RECT 5.3300 1.6550 5.5000 1.8700 ;
	    RECT 5.3300 1.2450 5.8950 1.6550 ;
	    RECT 5.3300 1.0300 5.5000 1.2450 ;
	    RECT 5.2150 0.8550 5.5000 1.0300 ;
	    RECT 5.2150 0.5200 5.4650 0.8550 ;
      END
   END Q
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 5.9800 3.5050 ;
	    RECT 0.5150 2.6700 0.8450 3.2950 ;
	    RECT 1.9750 2.2950 2.2900 3.2950 ;
	    RECT 3.8400 2.6700 4.1400 3.2950 ;
	    RECT 4.7600 1.8700 5.0450 3.2950 ;
	    RECT 5.6350 2.1950 5.8950 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.9800 3.7000 ;
      END
   END vpwr
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.8950 0.1050 2.2250 0.5550 ;
	    RECT 3.7600 0.1050 4.0900 1.0300 ;
	    RECT 4.7600 0.1050 5.0450 1.0300 ;
	    RECT 5.6350 0.1050 5.8950 0.6900 ;
	    RECT 0.0000 -0.1050 5.9800 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.9800 0.3000 ;
      END
   END vgnd
   OBS
         LAYER li1 ;
	    RECT 0.1750 2.4550 0.3450 3.0800 ;
	    RECT 0.1750 2.2450 0.7800 2.4550 ;
	    RECT 0.6100 1.7500 0.7800 2.2450 ;
	    RECT 1.0150 2.1050 1.2400 3.0800 ;
	    RECT 0.6100 1.3400 0.8400 1.7500 ;
	    RECT 0.6100 1.0050 0.7800 1.3400 ;
	    RECT 0.1750 0.7950 0.7800 1.0050 ;
	    RECT 0.1750 0.4300 0.3450 0.7950 ;
	    RECT 1.0150 0.4300 1.1850 2.1050 ;
	    RECT 1.4750 2.0800 1.8050 3.0200 ;
	    RECT 2.9200 2.8200 3.6700 3.0300 ;
	    RECT 1.4750 1.8700 2.1600 2.0800 ;
	    RECT 1.9900 1.3700 2.1600 1.8700 ;
	    RECT 2.4900 1.6950 2.7750 2.5050 ;
	    RECT 2.9450 1.7700 3.2850 2.4950 ;
	    RECT 1.9900 0.9800 2.3600 1.3700 ;
	    RECT 2.9450 1.2950 3.1150 1.7700 ;
	    RECT 3.5000 1.6550 3.6700 2.8200 ;
	    RECT 4.3600 2.3300 4.5800 3.0450 ;
	    RECT 3.8600 1.9200 4.5800 2.3300 ;
	    RECT 4.4100 1.6550 4.5800 1.9200 ;
	    RECT 3.5000 1.4550 4.2200 1.6550 ;
	    RECT 1.5550 0.9550 2.3600 0.9800 ;
	    RECT 1.5550 0.7700 2.1600 0.9550 ;
	    RECT 2.7350 0.8800 3.1150 1.2950 ;
	    RECT 3.3500 1.2450 4.2200 1.4550 ;
	    RECT 4.4100 1.2450 5.1600 1.6550 ;
	    RECT 1.5550 0.4300 1.7250 0.7700 ;
	    RECT 3.3500 0.6700 3.5200 1.2450 ;
	    RECT 4.4100 1.0300 4.5800 1.2450 ;
	    RECT 2.8600 0.4550 3.5200 0.6700 ;
	    RECT 4.3600 0.5200 4.5800 1.0300 ;
         LAYER met1 ;
	    RECT 1.0100 2.4250 1.3000 2.4800 ;
	    RECT 2.4300 2.4250 2.7200 2.4800 ;
	    RECT 1.0100 2.2500 2.7200 2.4250 ;
	    RECT 1.0100 2.1950 1.3000 2.2500 ;
	    RECT 2.4300 2.1950 2.7200 2.2500 ;
	    RECT 0.5500 2.0000 0.8400 2.0550 ;
	    RECT 2.8900 2.0000 3.1800 2.0550 ;
	    RECT 0.5500 1.8250 3.1800 2.0000 ;
	    RECT 0.5500 1.7700 0.8400 1.8250 ;
	    RECT 2.8900 1.7700 3.1800 1.8250 ;
   END
END efs8hd_dlxtn_2
MACRO efs8hd_dlygate4sd2_1
   CLASS CORE ;
   FOREIGN efs8hd_dlygate4sd2_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.2200 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 2.5700 1.8700 3.1350 3.0800 ;
	    RECT 2.6750 1.0300 3.1350 1.8700 ;
	    RECT 2.5700 0.3200 3.1350 1.0300 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3200 0.7750 2.0200 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.6550 0.1050 0.9250 0.6800 ;
	    RECT 2.0750 0.1050 2.4000 0.6800 ;
	    RECT 0.6550 0.0850 2.4000 0.1050 ;
	    RECT 0.0000 -0.0850 3.2200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.2200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.2200 3.4850 ;
	    RECT 0.6550 3.2950 2.4000 3.3150 ;
	    RECT 0.6550 2.7200 0.9250 3.2950 ;
	    RECT 2.0750 2.7200 2.4000 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.2200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.5050 0.4850 3.0800 ;
	    RECT 1.1550 2.6750 1.4550 3.0800 ;
	    RECT 0.0850 2.2300 1.1150 2.5050 ;
	    RECT 0.9450 1.1050 1.1150 2.2300 ;
	    RECT 0.0850 0.9000 1.1150 1.1050 ;
	    RECT 1.2850 2.0200 1.4550 2.6750 ;
	    RECT 1.6250 2.5050 1.8750 3.0800 ;
	    RECT 1.6250 2.2300 2.4000 2.5050 ;
	    RECT 1.2850 1.3200 2.0300 2.0200 ;
	    RECT 2.2000 1.6550 2.4000 2.2300 ;
	    RECT 0.0850 0.3200 0.4850 0.9000 ;
	    RECT 1.2850 0.7300 1.4550 1.3200 ;
	    RECT 2.2000 1.2450 2.5050 1.6550 ;
	    RECT 2.2000 1.1050 2.4000 1.2450 ;
	    RECT 1.1550 0.3200 1.4550 0.7300 ;
	    RECT 1.6250 0.8950 2.4000 1.1050 ;
	    RECT 1.6250 0.3200 1.8750 0.8950 ;
   END
END efs8hd_dlygate4sd2_1
MACRO efs8hd_dlygate4sd3_1
   CLASS CORE ;
   FOREIGN efs8hd_dlygate4sd3_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.6800 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3200 0.7750 2.0200 ;
      END
   END A
   PIN X
      PORT
         LAYER li1 ;
	    RECT 3.2100 1.8700 3.5950 3.0800 ;
	    RECT 3.3150 1.0300 3.5950 1.8700 ;
	    RECT 3.2100 0.3200 3.5950 1.0300 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.6550 0.1050 0.9250 0.6800 ;
	    RECT 2.7150 0.1050 3.0400 0.6800 ;
	    RECT 0.0000 -0.1050 3.6800 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.6800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 3.6800 3.5050 ;
	    RECT 0.6550 2.7200 0.9250 3.2950 ;
	    RECT 2.7150 2.7200 3.0400 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.6800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.2000 2.5050 0.4850 3.0800 ;
	    RECT 0.2000 2.2300 1.1550 2.5050 ;
	    RECT 0.9450 1.1050 1.1550 2.2300 ;
	    RECT 0.2000 0.8950 1.1550 1.1050 ;
	    RECT 1.3250 2.0200 1.7250 3.0800 ;
	    RECT 1.9150 2.5050 2.1950 3.0800 ;
	    RECT 1.9150 2.2300 3.0400 2.5050 ;
	    RECT 1.3250 1.3200 2.4200 2.0200 ;
	    RECT 2.5900 1.6550 3.0400 2.2300 ;
	    RECT 0.2000 0.3200 0.4850 0.8950 ;
	    RECT 1.3250 0.3200 1.7250 1.3200 ;
	    RECT 2.5900 1.2450 3.1450 1.6550 ;
	    RECT 2.5900 1.1050 3.0400 1.2450 ;
	    RECT 1.9150 0.8950 3.0400 1.1050 ;
	    RECT 1.9150 0.3200 2.1950 0.8950 ;
   END
END efs8hd_dlygate4sd3_1
MACRO efs8hd_dlymetal6s2s_1
   CLASS CORE ;
   FOREIGN efs8hd_dlymetal6s2s_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.6000 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 1.2450 2.0950 1.6700 3.0800 ;
	    RECT 1.2450 1.8700 2.1550 2.0950 ;
	    RECT 1.3200 1.2450 2.1550 1.8700 ;
	    RECT 1.3200 1.0300 1.6700 1.2450 ;
	    RECT 1.2450 0.3200 1.6700 1.0300 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.1050 0.5700 2.1250 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.6900 0.1050 1.0750 0.5950 ;
	    RECT 2.2850 0.1050 2.6700 0.6050 ;
	    RECT 3.7000 0.1050 4.0850 0.6050 ;
	    RECT 0.6900 0.0850 4.0850 0.1050 ;
	    RECT 0.0000 -0.0850 4.6000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.6000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.6000 3.4850 ;
	    RECT 0.6900 3.2950 4.0850 3.3150 ;
	    RECT 0.6900 2.7650 1.0750 3.2950 ;
	    RECT 2.2850 2.7650 2.6700 3.2950 ;
	    RECT 3.7000 2.7650 4.0850 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.6000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.5500 0.5200 3.0800 ;
	    RECT 1.8400 2.5500 2.1150 3.0800 ;
	    RECT 0.0850 2.3400 1.0750 2.5500 ;
	    RECT 0.7400 1.6550 1.0750 2.3400 ;
	    RECT 1.8400 2.3050 2.6700 2.5500 ;
	    RECT 2.3250 1.6550 2.6700 2.3050 ;
	    RECT 2.8400 2.0950 3.0850 3.0800 ;
	    RECT 3.2750 2.5500 3.5300 3.0800 ;
	    RECT 3.2750 2.3050 4.0850 2.5500 ;
	    RECT 2.8400 1.8700 3.5650 2.0950 ;
	    RECT 0.7400 1.2450 1.1500 1.6550 ;
	    RECT 2.3250 1.2450 2.7450 1.6550 ;
	    RECT 2.9150 1.2450 3.5650 1.8700 ;
	    RECT 3.7350 1.6550 4.0850 2.3050 ;
	    RECT 4.2550 1.8700 4.5150 3.0800 ;
	    RECT 3.7350 1.2450 4.1600 1.6550 ;
	    RECT 0.7400 0.9350 1.0750 1.2450 ;
	    RECT 2.3250 1.0300 2.6700 1.2450 ;
	    RECT 2.9150 1.0300 3.0850 1.2450 ;
	    RECT 3.7350 1.0300 4.0850 1.2450 ;
	    RECT 4.3300 1.0300 4.5150 1.8700 ;
	    RECT 0.0850 0.7650 1.0750 0.9350 ;
	    RECT 1.8600 0.8200 2.6700 1.0300 ;
	    RECT 0.0850 0.3200 0.5200 0.7650 ;
	    RECT 1.8600 0.3200 2.1150 0.8200 ;
	    RECT 2.8400 0.3200 3.0850 1.0300 ;
	    RECT 3.2750 0.8200 4.0850 1.0300 ;
	    RECT 3.2750 0.3200 3.5300 0.8200 ;
	    RECT 4.2550 0.3200 4.5150 1.0300 ;
   END
END efs8hd_dlymetal6s2s_1
MACRO efs8hd_dlymetal6s4s_1
   CLASS CORE ;
   FOREIGN efs8hd_dlymetal6s4s_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.6000 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 2.6600 2.0950 3.1050 3.0800 ;
	    RECT 2.6600 1.8700 3.5650 2.0950 ;
	    RECT 2.7350 1.2450 3.5650 1.8700 ;
	    RECT 2.7350 1.0300 3.1050 1.2450 ;
	    RECT 2.6600 0.3200 3.1050 1.0300 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.1050 0.5700 2.1250 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.6900 0.1050 1.0750 0.5950 ;
	    RECT 2.1050 0.1050 2.4900 0.6050 ;
	    RECT 3.7000 0.1050 4.0850 0.6050 ;
	    RECT 0.6900 0.0850 4.0850 0.1050 ;
	    RECT 0.0000 -0.0850 4.6000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.6000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.6000 3.4850 ;
	    RECT 0.6900 3.2950 4.0850 3.3150 ;
	    RECT 0.6900 2.7650 1.0750 3.2950 ;
	    RECT 2.1050 2.7650 2.4900 3.2950 ;
	    RECT 3.7000 2.7650 4.0850 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.6000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.5500 0.5200 3.0800 ;
	    RECT 0.0850 2.3400 1.0750 2.5500 ;
	    RECT 0.7400 1.6550 1.0750 2.3400 ;
	    RECT 1.2450 2.0950 1.5150 3.0800 ;
	    RECT 1.6850 2.5500 1.9350 3.0800 ;
	    RECT 3.2750 2.5500 3.5300 3.0800 ;
	    RECT 1.6850 2.3050 2.4900 2.5500 ;
	    RECT 3.2750 2.3050 4.0850 2.5500 ;
	    RECT 1.2450 1.8700 1.9700 2.0950 ;
	    RECT 0.7400 1.2450 1.1500 1.6550 ;
	    RECT 1.3200 1.2450 1.9700 1.8700 ;
	    RECT 2.1400 1.6550 2.4900 2.3050 ;
	    RECT 3.7350 1.6550 4.0850 2.3050 ;
	    RECT 4.2550 1.8700 4.5150 3.0800 ;
	    RECT 2.1400 1.2450 2.5650 1.6550 ;
	    RECT 3.7350 1.2450 4.1600 1.6550 ;
	    RECT 0.7400 0.9350 1.0750 1.2450 ;
	    RECT 1.3200 1.0300 1.5150 1.2450 ;
	    RECT 2.1400 1.0300 2.4900 1.2450 ;
	    RECT 3.7350 1.0300 4.0850 1.2450 ;
	    RECT 4.3300 1.0300 4.5150 1.8700 ;
	    RECT 0.0850 0.7650 1.0750 0.9350 ;
	    RECT 0.0850 0.3200 0.5200 0.7650 ;
	    RECT 1.2450 0.3200 1.5150 1.0300 ;
	    RECT 1.6850 0.8200 2.4900 1.0300 ;
	    RECT 3.2750 0.8200 4.0850 1.0300 ;
	    RECT 1.6850 0.3200 1.9350 0.8200 ;
	    RECT 3.2750 0.3200 3.5300 0.8200 ;
	    RECT 4.2550 0.3200 4.5150 1.0300 ;
   END
END efs8hd_dlymetal6s4s_1
MACRO efs8hd_dlymetal6s6s_1
   CLASS CORE ;
   FOREIGN efs8hd_dlymetal6s6s_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.6000 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 4.0800 1.8700 4.5150 3.0800 ;
	    RECT 4.1550 1.0300 4.5150 1.8700 ;
	    RECT 4.0800 0.3200 4.5150 1.0300 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.1050 0.5750 2.1250 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.6950 0.1050 1.0800 0.5950 ;
	    RECT 2.1100 0.1050 2.4950 0.6050 ;
	    RECT 3.5250 0.1050 3.9100 0.6050 ;
	    RECT 0.6950 0.0850 3.9100 0.1050 ;
	    RECT 0.0000 -0.0850 4.6000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.6000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.6000 3.4850 ;
	    RECT 0.6950 3.2950 3.9100 3.3150 ;
	    RECT 0.6950 2.7650 1.0800 3.2950 ;
	    RECT 2.1100 2.7650 2.4950 3.2950 ;
	    RECT 3.5250 2.7650 3.9100 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.6000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.5500 0.5250 3.0800 ;
	    RECT 0.0850 2.3400 1.0800 2.5500 ;
	    RECT 0.7450 1.6550 1.0800 2.3400 ;
	    RECT 1.2500 2.0950 1.5200 3.0800 ;
	    RECT 1.6900 2.5500 1.9400 3.0800 ;
	    RECT 1.6900 2.3050 2.4950 2.5500 ;
	    RECT 1.2500 1.8700 1.9750 2.0950 ;
	    RECT 0.7450 1.2450 1.1550 1.6550 ;
	    RECT 1.3250 1.2450 1.9750 1.8700 ;
	    RECT 2.1450 1.6550 2.4950 2.3050 ;
	    RECT 2.6650 2.0950 2.9150 3.0800 ;
	    RECT 3.0850 2.5500 3.3550 3.0800 ;
	    RECT 3.0850 2.3050 3.9100 2.5500 ;
	    RECT 2.6650 1.8700 3.3900 2.0950 ;
	    RECT 2.1450 1.2450 2.5700 1.6550 ;
	    RECT 2.7400 1.2450 3.3900 1.8700 ;
	    RECT 3.5600 1.6550 3.9100 2.3050 ;
	    RECT 3.5600 1.2450 3.9850 1.6550 ;
	    RECT 0.7450 0.9350 1.0800 1.2450 ;
	    RECT 1.3250 1.0300 1.5200 1.2450 ;
	    RECT 2.1450 1.0300 2.4950 1.2450 ;
	    RECT 2.7400 1.0300 2.9150 1.2450 ;
	    RECT 3.5600 1.0300 3.9100 1.2450 ;
	    RECT 0.0850 0.7650 1.0800 0.9350 ;
	    RECT 0.0850 0.3200 0.5250 0.7650 ;
	    RECT 1.2500 0.3200 1.5200 1.0300 ;
	    RECT 1.6900 0.8200 2.4950 1.0300 ;
	    RECT 1.6900 0.3200 1.9400 0.8200 ;
	    RECT 2.6650 0.3200 2.9150 1.0300 ;
	    RECT 3.0850 0.8200 3.9100 1.0300 ;
	    RECT 3.0850 0.3200 3.3550 0.8200 ;
   END
END efs8hd_dlymetal6s6s_1
MACRO efs8hd_einvn_1
   CLASS CORE ;
   FOREIGN efs8hd_einvn_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 2.8750 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 1.9700 0.9550 2.2150 2.0150 ;
      END
   END A
   PIN TEB
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.1900 0.5100 2.1550 ;
      END
   END TEB
   PIN Z
      PORT
         LAYER li1 ;
	    RECT 1.0400 2.2300 2.2150 3.0800 ;
	    RECT 1.6200 0.7400 1.8000 2.2300 ;
	    RECT 1.6200 0.3150 2.2150 0.7400 ;
      END
   END Z
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5400 0.0850 1.4400 0.5550 ;
	    RECT 0.0000 -0.0850 2.3000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 2.3000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 2.3000 3.4850 ;
	    RECT 0.5400 2.7900 0.8700 3.3150 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 2.3000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.5800 0.3700 3.0800 ;
	    RECT 0.0850 2.3650 0.8700 2.5800 ;
	    RECT 0.6850 2.0150 0.8700 2.3650 ;
	    RECT 0.6850 0.9800 1.4500 2.0150 ;
	    RECT 0.0850 0.7650 1.4500 0.9800 ;
	    RECT 0.0850 0.3150 0.3700 0.7650 ;
   END
END efs8hd_einvn_1
MACRO efs8hd_einvn_2
   CLASS CORE ;
   FOREIGN efs8hd_einvn_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.0250 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 2.7850 1.3400 3.1350 1.5900 ;
      END
   END A
   PIN TEB
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.2400 0.3250 1.7300 ;
      END
   END TEB
   PIN Z
      PORT
         LAYER li1 ;
	    RECT 2.7850 2.1150 3.1350 3.0800 ;
	    RECT 1.9450 1.8050 3.1350 2.1150 ;
	    RECT 2.3650 1.0550 2.6150 1.8050 ;
	    RECT 2.3650 0.7400 2.6950 1.0550 ;
      END
   END Z
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.0850 0.8450 0.6050 ;
	    RECT 1.4500 0.0850 1.7800 0.6050 ;
	    RECT 0.0000 -0.0850 3.2200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.2200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.2200 3.4850 ;
	    RECT 0.5150 2.3650 0.8950 3.3150 ;
	    RECT 1.4100 2.8150 2.2750 3.3150 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.2200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.1550 0.3450 3.0800 ;
	    RECT 1.0700 2.6050 1.2400 3.0800 ;
	    RECT 2.4450 2.6050 2.6150 3.0800 ;
	    RECT 1.0700 2.3300 2.6150 2.6050 ;
	    RECT 0.0850 1.9400 0.8950 2.1550 ;
	    RECT 0.4950 1.5900 0.8950 1.9400 ;
	    RECT 1.0700 1.8050 1.7750 2.3300 ;
	    RECT 0.4950 1.2400 2.0350 1.5900 ;
	    RECT 0.4950 1.0300 0.8400 1.2400 ;
	    RECT 0.0850 0.8150 0.8400 1.0300 ;
	    RECT 1.0150 0.8150 2.1950 1.0300 ;
	    RECT 0.0850 0.3150 0.3450 0.8150 ;
	    RECT 1.0150 0.3150 1.2800 0.8150 ;
	    RECT 1.9500 0.5300 2.1950 0.8150 ;
	    RECT 2.8650 0.5300 3.1350 0.9650 ;
	    RECT 1.9500 0.3150 3.1350 0.5300 ;
   END
END efs8hd_einvn_2
MACRO efs8hd_einvn_4
   CLASS CORE ;
   FOREIGN efs8hd_einvn_4 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 6.3250 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 4.5300 0.7750 4.9750 1.6550 ;
      END
   END A
   PIN TEB
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.2400 0.3450 1.6550 ;
      END
   END TEB
   PIN Z
      PORT
         LAYER li1 ;
	    RECT 3.1900 1.8500 3.5200 2.5900 ;
	    RECT 4.0300 1.8500 4.3600 2.5900 ;
	    RECT 3.1900 0.7750 4.3600 1.8500 ;
      END
   END Z
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.0850 0.8450 0.6050 ;
	    RECT 1.4550 0.0850 1.7850 0.6050 ;
	    RECT 2.2950 0.0850 2.6250 0.6050 ;
	    RECT 0.0000 -0.0850 5.0600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.0600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.0600 3.4850 ;
	    RECT 0.5150 2.2900 0.8450 3.3150 ;
	    RECT 1.4100 2.2900 1.7400 3.3150 ;
	    RECT 2.2500 2.2900 2.6400 3.3150 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.0600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.0800 0.3450 3.0800 ;
	    RECT 1.0150 2.0800 1.2400 3.0800 ;
	    RECT 1.9100 2.0800 2.0800 3.0800 ;
	    RECT 2.8100 2.8650 4.9750 3.0800 ;
	    RECT 2.8100 2.0800 3.0200 2.8650 ;
	    RECT 0.0850 1.8650 0.8450 2.0800 ;
	    RECT 1.0150 1.8650 3.0200 2.0800 ;
	    RECT 3.6900 2.0600 3.8600 2.8650 ;
	    RECT 4.5300 2.0600 4.9750 2.8650 ;
	    RECT 0.5150 1.6550 0.8450 1.8650 ;
	    RECT 0.5150 1.2400 3.0200 1.6550 ;
	    RECT 0.5150 1.0300 0.8450 1.2400 ;
	    RECT 0.0850 0.8150 0.8450 1.0300 ;
	    RECT 1.0150 0.8150 2.9950 1.0300 ;
	    RECT 0.0850 0.3150 0.3450 0.8150 ;
	    RECT 1.0150 0.3150 1.2850 0.8150 ;
	    RECT 1.9550 0.3150 2.1250 0.8150 ;
	    RECT 2.8250 0.5600 2.9950 0.8150 ;
	    RECT 2.8250 0.3150 4.9750 0.5600 ;
   END
END efs8hd_einvn_4
MACRO efs8hd_einvn_8
   CLASS CORE ;
   FOREIGN efs8hd_einvn_8 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 10.3500 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 4.6450 1.2400 7.8000 1.6050 ;
      END
   END A
   PIN TEB
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.2400 0.3450 1.6550 ;
      END
   END TEB
   PIN Z
      PORT
         LAYER li1 ;
	    RECT 4.8700 2.0300 5.2000 2.6550 ;
	    RECT 5.7100 2.0300 6.0400 2.6550 ;
	    RECT 6.5500 2.0300 6.8800 2.6550 ;
	    RECT 7.3900 2.0300 7.7200 2.6550 ;
	    RECT 4.8700 1.8150 8.1950 2.0300 ;
	    RECT 7.9700 1.0300 8.1950 1.8150 ;
	    RECT 4.8700 0.7750 8.1950 1.0300 ;
      END
   END Z
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.0850 0.8450 0.6050 ;
	    RECT 1.4550 0.0850 1.7850 0.6050 ;
	    RECT 2.2950 0.0850 2.6250 0.6050 ;
	    RECT 3.1350 0.0850 3.4650 0.6050 ;
	    RECT 3.9750 0.0850 4.3150 0.6050 ;
	    RECT 0.0000 -0.0850 8.2800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 8.2800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 8.2800 3.4850 ;
	    RECT 0.5150 2.2900 0.8450 3.3150 ;
	    RECT 1.4100 2.2900 1.7400 3.3150 ;
	    RECT 2.2500 2.2900 2.5800 3.3150 ;
	    RECT 3.0900 2.2900 3.4200 3.3150 ;
	    RECT 3.9300 2.2900 4.2800 3.3150 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 8.2800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0900 2.0800 0.3450 3.0800 ;
	    RECT 1.0150 2.0800 1.2400 3.0800 ;
	    RECT 1.9100 2.0800 2.0800 3.0800 ;
	    RECT 2.7500 2.0800 2.9200 3.0800 ;
	    RECT 3.5900 2.0800 3.7600 3.0800 ;
	    RECT 4.4500 2.8650 8.1950 3.0800 ;
	    RECT 4.4500 2.0800 4.7000 2.8650 ;
	    RECT 5.3700 2.2400 5.5400 2.8650 ;
	    RECT 6.2100 2.2400 6.3800 2.8650 ;
	    RECT 7.0500 2.2400 7.2200 2.8650 ;
	    RECT 7.8900 2.2400 8.1950 2.8650 ;
	    RECT 0.0900 1.8650 0.8450 2.0800 ;
	    RECT 1.0150 1.8650 4.7000 2.0800 ;
	    RECT 0.5150 1.6550 0.8450 1.8650 ;
	    RECT 0.5150 1.2400 4.4750 1.6550 ;
	    RECT 0.5150 1.0300 0.8450 1.2400 ;
	    RECT 0.0900 0.8150 0.8450 1.0300 ;
	    RECT 1.0150 0.8150 4.7000 1.0300 ;
	    RECT 0.0900 0.3150 0.3450 0.8150 ;
	    RECT 1.0150 0.3150 1.2850 0.8150 ;
	    RECT 1.9550 0.3150 2.1250 0.8150 ;
	    RECT 2.7950 0.3150 2.9650 0.8150 ;
	    RECT 3.6350 0.3150 3.8050 0.8150 ;
	    RECT 4.4850 0.5600 4.7000 0.8150 ;
	    RECT 4.4850 0.3150 8.1950 0.5600 ;
   END
END efs8hd_einvn_8
MACRO efs8hd_einvp_1
   CLASS CORE ;
   FOREIGN efs8hd_einvp_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 2.8750 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 1.9750 1.2150 2.2150 2.4400 ;
      END
   END A
   PIN TE
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.2400 0.5450 2.1550 ;
      END
   END TE
   PIN Z
      PORT
         LAYER li1 ;
	    RECT 1.6200 2.6550 2.2150 3.0800 ;
	    RECT 1.6200 1.0050 1.7950 2.6550 ;
	    RECT 1.6200 0.3150 2.2150 1.0050 ;
      END
   END Z
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.0850 1.4500 0.6050 ;
	    RECT 0.0000 -0.0850 2.3000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 2.3000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 2.3000 3.4850 ;
	    RECT 0.5150 2.7900 1.4500 3.3150 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 2.3000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.5800 0.3450 3.0800 ;
	    RECT 0.0850 2.3650 1.4500 2.5800 ;
	    RECT 0.7150 1.0300 1.4500 2.3650 ;
	    RECT 0.0850 0.8150 1.4500 1.0300 ;
	    RECT 0.0850 0.3150 0.3450 0.8150 ;
   END
END efs8hd_einvp_1
MACRO efs8hd_einvp_2
   CLASS CORE ;
   FOREIGN efs8hd_einvp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.0250 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 2.8500 0.9550 3.1350 2.0150 ;
      END
   END A
   PIN TE
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.2400 0.3300 2.0150 ;
      END
   END TE
   PIN Z
      PORT
         LAYER li1 ;
	    RECT 2.3500 0.7400 2.6800 2.6550 ;
      END
   END Z
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.0850 0.8750 0.6050 ;
	    RECT 1.4100 0.0850 1.7700 0.6050 ;
	    RECT 0.0000 -0.0850 3.2200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.2200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.2200 3.4850 ;
	    RECT 0.5150 2.6550 0.8750 3.3150 ;
	    RECT 1.4550 2.3650 1.7850 3.3150 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.2200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.4400 0.3450 3.0800 ;
	    RECT 0.0850 2.2300 0.8750 2.4400 ;
	    RECT 0.5000 1.6550 0.8750 2.2300 ;
	    RECT 1.0450 2.1550 1.2850 3.0800 ;
	    RECT 1.9850 2.8650 3.1350 3.0800 ;
	    RECT 1.9850 2.1550 2.1550 2.8650 ;
	    RECT 2.8500 2.2300 3.1350 2.8650 ;
	    RECT 1.0450 1.9400 2.1550 2.1550 ;
	    RECT 0.5000 1.2400 2.1800 1.6550 ;
	    RECT 0.5000 1.0300 0.8750 1.2400 ;
	    RECT 0.0850 0.8150 0.8750 1.0300 ;
	    RECT 1.0450 0.8150 2.1800 1.0300 ;
	    RECT 0.0850 0.3150 0.3450 0.8150 ;
	    RECT 1.0450 0.3150 1.2400 0.8150 ;
	    RECT 1.9400 0.5300 2.1800 0.8150 ;
	    RECT 2.8500 0.5300 3.1350 0.7400 ;
	    RECT 1.9400 0.3150 3.1350 0.5300 ;
   END
END efs8hd_einvp_2
MACRO efs8hd_einvp_4
   CLASS CORE ;
   FOREIGN efs8hd_einvp_4 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 6.3250 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 3.7400 1.2750 4.9750 1.5900 ;
      END
   END A
   PIN TE
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.2400 0.3300 2.0150 ;
      END
   END TE
   PIN Z
      PORT
         LAYER li1 ;
	    RECT 3.1900 2.0150 3.5200 2.6550 ;
	    RECT 4.0300 2.0150 4.3600 2.6550 ;
	    RECT 3.1900 1.8050 4.3600 2.0150 ;
	    RECT 3.1900 1.0600 3.5700 1.8050 ;
	    RECT 3.1900 0.7900 4.9750 1.0600 ;
      END
   END Z
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.0850 0.8450 0.6050 ;
	    RECT 1.3750 0.0850 1.7050 0.6050 ;
	    RECT 2.2150 0.0850 2.5550 0.6050 ;
	    RECT 0.0000 -0.0850 5.0600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.0600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.0600 3.4850 ;
	    RECT 0.5150 2.6550 0.8750 3.3150 ;
	    RECT 1.4550 2.3650 1.7850 3.3150 ;
	    RECT 2.2950 2.3650 2.6550 3.3150 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.0600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.4400 0.3450 3.0800 ;
	    RECT 0.0850 2.2300 0.8750 2.4400 ;
	    RECT 0.5000 1.6550 0.8750 2.2300 ;
	    RECT 1.0750 2.1550 1.2850 3.0800 ;
	    RECT 1.9550 2.1550 2.1250 3.0800 ;
	    RECT 2.8250 2.8650 4.9750 3.0800 ;
	    RECT 2.8250 2.1550 2.9950 2.8650 ;
	    RECT 3.6900 2.2300 3.8600 2.8650 ;
	    RECT 1.0750 1.9400 2.9950 2.1550 ;
	    RECT 4.5300 1.8050 4.9750 2.8650 ;
	    RECT 0.5000 1.2400 3.0200 1.6550 ;
	    RECT 0.5000 1.0300 0.6950 1.2400 ;
	    RECT 0.0850 0.8150 0.6950 1.0300 ;
	    RECT 1.0350 0.8150 3.0200 1.0300 ;
	    RECT 0.0850 0.3150 0.3450 0.8150 ;
	    RECT 1.0350 0.3150 1.2050 0.8150 ;
	    RECT 1.8750 0.3150 2.0450 0.8150 ;
	    RECT 2.7350 0.5800 3.0200 0.8150 ;
	    RECT 2.7350 0.3150 4.9750 0.5800 ;
   END
END efs8hd_einvp_4
MACRO efs8hd_einvp_8
   CLASS CORE ;
   FOREIGN efs8hd_einvp_8 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 10.3500 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 5.4200 1.2750 8.1950 1.5900 ;
      END
   END A
   PIN TE
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.2400 0.3300 2.0150 ;
      END
   END TE
   PIN Z
      PORT
         LAYER li1 ;
	    RECT 4.8700 2.0150 5.2000 2.6550 ;
	    RECT 5.7100 2.0150 6.0400 2.6550 ;
	    RECT 6.5500 2.0150 6.8800 2.6550 ;
	    RECT 7.3900 2.0150 7.7200 2.6550 ;
	    RECT 4.8700 1.8050 7.7200 2.0150 ;
	    RECT 4.8700 1.0600 5.2500 1.8050 ;
	    RECT 4.8700 0.7900 8.1950 1.0600 ;
      END
   END Z
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.0850 0.8450 0.6050 ;
	    RECT 1.3750 0.0850 1.7050 0.6050 ;
	    RECT 2.2150 0.0850 2.5450 0.6050 ;
	    RECT 3.0550 0.0850 3.3850 0.6050 ;
	    RECT 3.8950 0.0850 4.2350 0.6050 ;
	    RECT 0.0000 -0.0850 8.2800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 8.2800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 8.2800 3.4850 ;
	    RECT 0.5150 2.6550 0.8750 3.3150 ;
	    RECT 1.4550 2.3650 1.7850 3.3150 ;
	    RECT 2.2950 2.3650 2.6250 3.3150 ;
	    RECT 3.1350 2.3650 3.4650 3.3150 ;
	    RECT 3.9750 2.3650 4.3050 3.3150 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 8.2800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.4400 0.3450 3.0800 ;
	    RECT 0.0850 2.2300 0.8750 2.4400 ;
	    RECT 0.5000 1.6550 0.8750 2.2300 ;
	    RECT 1.0750 2.1550 1.2850 3.0800 ;
	    RECT 1.9550 2.1550 2.1250 3.0800 ;
	    RECT 2.7950 2.1550 2.9650 3.0800 ;
	    RECT 3.6350 2.1550 3.8050 3.0800 ;
	    RECT 4.4750 2.8650 8.1950 3.0800 ;
	    RECT 4.4750 2.1550 4.7000 2.8650 ;
	    RECT 5.3700 2.2300 5.5400 2.8650 ;
	    RECT 6.2100 2.2300 6.3800 2.8650 ;
	    RECT 7.0500 2.2300 7.2200 2.8650 ;
	    RECT 1.0750 1.9400 4.7000 2.1550 ;
	    RECT 7.8900 1.8050 8.1950 2.8650 ;
	    RECT 0.5000 1.2400 4.7000 1.6550 ;
	    RECT 0.5000 1.0300 0.6950 1.2400 ;
	    RECT 0.0850 0.8150 0.6950 1.0300 ;
	    RECT 1.0350 0.8150 4.7000 1.0300 ;
	    RECT 0.0850 0.3150 0.3450 0.8150 ;
	    RECT 1.0350 0.3150 1.2050 0.8150 ;
	    RECT 1.8750 0.3150 2.0450 0.8150 ;
	    RECT 2.7150 0.3150 2.8850 0.8150 ;
	    RECT 3.5550 0.3150 3.7250 0.8150 ;
	    RECT 4.4050 0.5800 4.7000 0.8150 ;
	    RECT 4.4050 0.3150 8.1950 0.5800 ;
   END
END efs8hd_einvp_8
MACRO efs8hd_fill_1
   CLASS CORE ;
   FOREIGN efs8hd_fill_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 0.4600 BY 3.4000 ;
   SITE unitehd ;
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 0.4600 3.4850 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 0.4600 3.7000 ;
      END
   END vpwr
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0000 -0.0850 0.4600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 0.4600 0.3000 ;
      END
   END vgnd
END efs8hd_fill_1
MACRO efs8hd_fill_2
   CLASS CORE ;
   FOREIGN efs8hd_fill_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 0.9200 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0000 -0.0850 0.9200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 0.9200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 0.9200 3.4850 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 0.9200 3.7000 ;
      END
   END vpwr
END efs8hd_fill_2
MACRO efs8hd_fill_4
   CLASS CORE ;
   FOREIGN efs8hd_fill_4 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 1.8400 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0000 -0.0850 1.8400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 1.8400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 1.8400 3.4850 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 1.8400 3.7000 ;
      END
   END vpwr
END efs8hd_fill_4
MACRO efs8hd_fill_8
   CLASS CORE ;
   FOREIGN efs8hd_fill_8 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.6800 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0000 -0.0850 3.6800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.6800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.6800 3.4850 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.6800 3.7000 ;
      END
   END vpwr
END efs8hd_fill_8
MACRO efs8hd_inv_12
   CLASS CORE ;
   FOREIGN efs8hd_inv_12 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.9800 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.6800 2.0800 1.0100 3.0800 ;
	    RECT 1.5200 2.0800 1.8500 3.0800 ;
	    RECT 2.3600 2.0800 2.6900 3.0800 ;
	    RECT 3.2000 2.0800 3.5300 3.0800 ;
	    RECT 4.0400 2.0800 4.3700 3.0800 ;
	    RECT 4.8800 2.0800 5.2100 3.0800 ;
	    RECT 0.0850 1.8700 5.8950 2.0800 ;
	    RECT 0.0850 1.1300 0.5100 1.8700 ;
	    RECT 5.5450 1.1300 5.8950 1.8700 ;
	    RECT 0.0850 0.8950 5.8950 1.1300 ;
	    RECT 0.6800 0.3200 1.0100 0.8950 ;
	    RECT 1.5200 0.3200 1.8500 0.8950 ;
	    RECT 2.3600 0.3200 2.6900 0.8950 ;
	    RECT 3.2000 0.3200 3.5300 0.8950 ;
	    RECT 4.0400 0.3200 4.3700 0.8950 ;
	    RECT 4.8800 0.3200 5.2100 0.8950 ;
      END
   END Y
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.6800 1.3450 5.2700 1.6550 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.2550 0.1050 0.5100 0.6800 ;
	    RECT 1.1800 0.1050 1.3500 0.6800 ;
	    RECT 2.0200 0.1050 2.1900 0.6800 ;
	    RECT 2.8600 0.1050 3.0300 0.6800 ;
	    RECT 3.7000 0.1050 3.8700 0.6800 ;
	    RECT 4.5400 0.1050 4.7100 0.6800 ;
	    RECT 5.5550 0.1050 5.8950 0.6800 ;
	    RECT 0.2550 0.0850 5.8950 0.1050 ;
	    RECT 0.0000 -0.0850 5.9800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.9800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.9800 3.4850 ;
	    RECT 0.2550 3.2950 5.8950 3.3150 ;
	    RECT 0.2550 2.2950 0.5100 3.2950 ;
	    RECT 1.1800 2.2950 1.3500 3.2950 ;
	    RECT 2.0200 2.2950 2.1900 3.2950 ;
	    RECT 2.8600 2.2950 3.0300 3.2950 ;
	    RECT 3.7000 2.2950 3.8700 3.2950 ;
	    RECT 4.5400 2.2950 4.7100 3.2950 ;
	    RECT 5.5550 2.2950 5.8950 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.9800 3.7000 ;
      END
   END vpwr
END efs8hd_inv_12
MACRO efs8hd_inv_16
   CLASS CORE ;
   FOREIGN efs8hd_inv_16 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 7.3600 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5800 2.0800 0.9100 3.0800 ;
	    RECT 1.4200 2.0800 1.7500 3.0800 ;
	    RECT 2.2600 2.0800 2.5900 3.0800 ;
	    RECT 3.1000 2.0800 3.4300 3.0800 ;
	    RECT 3.9400 2.0800 4.2700 3.0800 ;
	    RECT 4.7800 2.0800 5.1100 3.0800 ;
	    RECT 5.6200 2.0800 5.9500 3.0800 ;
	    RECT 6.4600 2.0800 6.7900 3.0800 ;
	    RECT 0.5800 1.8700 6.7900 2.0800 ;
	    RECT 6.4600 1.1300 6.7900 1.8700 ;
	    RECT 0.5800 0.8950 6.7900 1.1300 ;
	    RECT 0.5800 0.3200 0.9100 0.8950 ;
	    RECT 1.4200 0.3200 1.7500 0.8950 ;
	    RECT 2.2600 0.3200 2.5900 0.8950 ;
	    RECT 3.1000 0.3200 3.4300 0.8950 ;
	    RECT 3.9400 0.3200 4.2700 0.8950 ;
	    RECT 4.7800 0.3200 5.1100 0.8950 ;
	    RECT 5.6200 0.3200 5.9500 0.8950 ;
	    RECT 6.4600 0.3200 6.7900 0.8950 ;
      END
   END Y
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3450 5.5250 1.6450 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1800 0.1050 0.4100 1.1050 ;
	    RECT 1.0800 0.1050 1.2500 0.6800 ;
	    RECT 1.9200 0.1050 2.0900 0.6800 ;
	    RECT 2.7600 0.1050 2.9300 0.6800 ;
	    RECT 3.6000 0.1050 3.7700 0.6800 ;
	    RECT 4.4400 0.1050 4.6100 0.6800 ;
	    RECT 5.2800 0.1050 5.4500 0.6800 ;
	    RECT 6.1200 0.1050 6.2900 0.6800 ;
	    RECT 6.9600 0.1050 7.1700 1.1050 ;
	    RECT 0.1800 0.0850 7.1700 0.1050 ;
	    RECT 0.0000 -0.0850 7.3600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 7.3600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 7.3600 3.4850 ;
	    RECT 0.2000 3.2950 7.1700 3.3150 ;
	    RECT 0.2000 1.8550 0.4100 3.2950 ;
	    RECT 1.0800 2.2950 1.2500 3.2950 ;
	    RECT 1.9200 2.2950 2.0900 3.2950 ;
	    RECT 2.7600 2.2950 2.9300 3.2950 ;
	    RECT 3.6000 2.2950 3.7700 3.2950 ;
	    RECT 4.4400 2.2950 4.6100 3.2950 ;
	    RECT 5.2800 2.2950 5.4500 3.2950 ;
	    RECT 6.1200 2.2950 6.2900 3.2950 ;
	    RECT 6.9600 2.2950 7.1700 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 7.3600 3.7000 ;
      END
   END vpwr
END efs8hd_inv_16
MACRO efs8hd_inv_2
   CLASS CORE ;
   FOREIGN efs8hd_inv_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 1.3800 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5250 1.8550 0.8550 3.0800 ;
	    RECT 0.6050 1.1050 0.8550 1.8550 ;
	    RECT 0.5250 0.3200 0.8550 1.1050 ;
      END
   END Y
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.1050 1.3450 0.4350 1.6550 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1250 0.1050 0.3550 1.1300 ;
	    RECT 1.0250 0.1050 1.2350 1.1300 ;
	    RECT 0.1250 0.0850 1.2350 0.1050 ;
	    RECT 0.0000 -0.0850 1.3800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 1.3800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 1.3800 3.4850 ;
	    RECT 0.1250 3.2950 1.2350 3.3150 ;
	    RECT 0.1250 1.8700 0.3550 3.2950 ;
	    RECT 1.0250 1.8700 1.2350 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 1.3800 3.7000 ;
      END
   END vpwr
END efs8hd_inv_2
MACRO efs8hd_inv_4
   CLASS CORE ;
   FOREIGN efs8hd_inv_4 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 2.3000 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5650 2.0800 0.8950 3.0800 ;
	    RECT 1.4050 2.1050 1.7350 3.0800 ;
	    RECT 1.4050 2.0800 2.1700 2.1050 ;
	    RECT 0.5650 1.8700 2.1700 2.0800 ;
	    RECT 1.9050 1.1300 2.1700 1.8700 ;
	    RECT 0.5650 0.9050 2.1700 1.1300 ;
	    RECT 0.5650 0.3200 0.8950 0.9050 ;
	    RECT 1.4050 0.3200 1.7350 0.9050 ;
      END
   END Y
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.1050 1.3450 1.7350 1.6550 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1300 0.1050 0.3950 0.6800 ;
	    RECT 1.0650 0.1050 1.2350 0.6800 ;
	    RECT 1.9050 0.1050 2.1550 0.6900 ;
	    RECT 0.1300 0.0850 2.1550 0.1050 ;
	    RECT 0.0000 -0.0850 2.3000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 2.3000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 2.3000 3.4850 ;
	    RECT 0.1300 3.2950 2.1150 3.3150 ;
	    RECT 0.1300 1.8700 0.3950 3.2950 ;
	    RECT 1.0650 2.2950 1.2350 3.2950 ;
	    RECT 1.9050 2.7200 2.1150 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 2.3000 3.7000 ;
      END
   END vpwr
END efs8hd_inv_4
MACRO efs8hd_inv_6
   CLASS CORE ;
   FOREIGN efs8hd_inv_6 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.2200 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.6850 2.0800 1.0150 3.0800 ;
	    RECT 1.5250 2.0800 1.8550 3.0800 ;
	    RECT 2.3650 2.1050 2.6950 3.0800 ;
	    RECT 2.3650 2.0800 3.1350 2.1050 ;
	    RECT 0.6850 1.8700 3.1350 2.0800 ;
	    RECT 2.7850 1.1300 3.1350 1.8700 ;
	    RECT 0.7650 0.9050 3.1350 1.1300 ;
	    RECT 0.7650 0.3200 0.9350 0.9050 ;
	    RECT 1.6050 0.3200 1.7750 0.9050 ;
	    RECT 2.4450 0.3200 2.6150 0.9050 ;
      END
   END Y
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.1050 1.3450 2.6150 1.6550 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1300 0.1050 0.3950 0.6800 ;
	    RECT 1.1850 0.1050 1.3550 0.6800 ;
	    RECT 2.0250 0.1050 2.1950 0.6800 ;
	    RECT 2.7850 0.1050 3.0350 0.6900 ;
	    RECT 0.1300 0.0850 3.0350 0.1050 ;
	    RECT 0.0000 -0.0850 3.2200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.2200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.2200 3.4850 ;
	    RECT 0.1300 3.2950 3.0350 3.3150 ;
	    RECT 0.1300 1.8700 0.4250 3.2950 ;
	    RECT 1.1850 2.2950 1.3550 3.2950 ;
	    RECT 2.0250 2.2950 2.1950 3.2950 ;
	    RECT 2.8650 2.7200 3.0350 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.2200 3.7000 ;
      END
   END vpwr
END efs8hd_inv_6
MACRO efs8hd_inv_8
   CLASS CORE ;
   FOREIGN efs8hd_inv_8 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.1400 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.6800 2.0800 1.0100 3.0800 ;
	    RECT 1.5200 2.0800 1.8500 3.0800 ;
	    RECT 2.3600 2.0800 2.6900 3.0800 ;
	    RECT 3.2000 2.0800 3.5300 3.0800 ;
	    RECT 0.0850 1.8700 4.0550 2.0800 ;
	    RECT 0.0850 1.1300 0.4300 1.8700 ;
	    RECT 3.7350 1.1300 4.0550 1.8700 ;
	    RECT 0.0850 0.8950 4.0550 1.1300 ;
	    RECT 0.6800 0.3200 1.0100 0.8950 ;
	    RECT 1.5200 0.3200 1.8500 0.8950 ;
	    RECT 2.3600 0.3200 2.6900 0.8950 ;
	    RECT 3.2000 0.3200 3.5300 0.8950 ;
      END
   END Y
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.6800 1.3450 3.5350 1.6550 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.2550 0.1050 0.5100 0.6800 ;
	    RECT 1.1800 0.1050 1.3500 0.6800 ;
	    RECT 2.0200 0.1050 2.1900 0.6800 ;
	    RECT 2.8600 0.1050 3.0300 0.6800 ;
	    RECT 3.7000 0.1050 4.0050 0.6800 ;
	    RECT 0.2550 0.0850 4.0050 0.1050 ;
	    RECT 0.0000 -0.0850 4.1400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.1400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.1400 3.4850 ;
	    RECT 0.2550 3.2950 4.0000 3.3150 ;
	    RECT 0.2550 2.2950 0.5100 3.2950 ;
	    RECT 1.1800 2.2950 1.3500 3.2950 ;
	    RECT 2.0200 2.2950 2.1900 3.2950 ;
	    RECT 2.8600 2.2950 3.0300 3.2950 ;
	    RECT 3.7000 2.2950 4.0000 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.1400 3.7000 ;
      END
   END vpwr
END efs8hd_inv_8
MACRO efs8hd_nand2_2
   CLASS CORE ;
   FOREIGN efs8hd_nand2_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 2.3000 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5150 2.0800 0.8450 3.0800 ;
	    RECT 1.3550 2.0800 1.6850 3.0800 ;
	    RECT 0.5150 1.8700 2.2150 2.0800 ;
	    RECT 1.9350 1.1300 2.2150 1.8700 ;
	    RECT 1.3550 0.8200 2.2150 1.1300 ;
      END
   END Y
   PIN B
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3450 0.8450 1.6550 ;
      END
   END B
   PIN A
      PORT
         LAYER li1 ;
	    RECT 1.0150 1.3450 1.7650 1.6550 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5950 0.0850 0.7650 0.6800 ;
	    RECT 0.0000 -0.0850 2.3000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 2.3000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 2.3000 3.4850 ;
	    RECT 0.0850 3.2950 2.1100 3.3150 ;
	    RECT 0.0850 1.8700 0.3450 3.2950 ;
	    RECT 1.0150 2.2950 1.1850 3.2950 ;
	    RECT 1.8550 2.2950 2.1100 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 2.3000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 0.8950 1.1850 1.1050 ;
	    RECT 0.0850 0.3200 0.4250 0.8950 ;
	    RECT 0.9350 0.5800 1.1850 0.8950 ;
	    RECT 1.7750 0.5800 2.1050 0.6050 ;
	    RECT 0.9350 0.3200 2.1050 0.5800 ;
   END
END efs8hd_nand2_2
MACRO efs8hd_nand2b_2
   CLASS CORE ;
   FOREIGN efs8hd_nand2b_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.2200 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 1.0350 2.5050 1.3650 3.0800 ;
	    RECT 2.2800 2.5050 2.6350 3.0800 ;
	    RECT 1.0350 2.2950 2.6350 2.5050 ;
	    RECT 1.5300 1.1300 1.8100 2.2950 ;
	    RECT 2.3600 1.8700 2.6350 2.2950 ;
	    RECT 1.5300 1.0050 1.8550 1.1300 ;
	    RECT 1.5250 0.7950 1.8550 1.0050 ;
      END
   END Y
   PIN AN
      PORT
         LAYER li1 ;
	    RECT 0.4550 1.1050 0.8000 1.6550 ;
      END
   END AN
   PIN B
      PORT
         LAYER li1 ;
	    RECT 1.9850 1.6150 2.1800 2.0700 ;
	    RECT 1.9850 1.3450 3.1350 1.6150 ;
      END
   END B
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.9350 ;
	    RECT 2.4450 0.1050 2.6150 0.6550 ;
	    RECT 0.5150 0.0850 2.6150 0.1050 ;
	    RECT 0.0000 -0.0850 3.2200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.2200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.2200 3.4850 ;
	    RECT 0.5800 3.2950 3.1350 3.3150 ;
	    RECT 0.5800 2.2950 0.8350 3.2950 ;
	    RECT 1.5350 2.7200 2.1100 3.2950 ;
	    RECT 2.8050 1.8700 3.1350 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.2200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1100 2.0800 0.4100 2.3250 ;
	    RECT 0.1100 1.8700 1.3600 2.0800 ;
	    RECT 0.1100 0.9750 0.2800 1.8700 ;
	    RECT 1.0300 1.3450 1.3600 1.8700 ;
	    RECT 0.1100 0.6400 0.3450 0.9750 ;
	    RECT 1.0800 0.5800 1.3550 1.1300 ;
	    RECT 2.0250 0.8700 3.1350 1.1300 ;
	    RECT 2.0250 0.5800 2.2750 0.8700 ;
	    RECT 1.0800 0.3200 2.2750 0.5800 ;
	    RECT 2.7850 0.3200 3.1350 0.8700 ;
   END
END efs8hd_nand2b_2
MACRO efs8hd_nand3_2
   CLASS CORE ;
   FOREIGN efs8hd_nand3_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.6800 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5150 2.0800 0.8450 3.0800 ;
	    RECT 1.3550 2.0800 1.6850 3.0800 ;
	    RECT 2.7150 2.0800 3.0450 3.0800 ;
	    RECT 0.5150 1.8050 3.0450 2.0800 ;
	    RECT 0.5150 0.7950 0.8450 1.8050 ;
      END
   END Y
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.1050 0.3300 1.6550 ;
      END
   END A
   PIN B
      PORT
         LAYER li1 ;
	    RECT 1.0650 1.3450 2.1600 1.6150 ;
      END
   END B
   PIN C
      PORT
         LAYER li1 ;
	    RECT 2.4450 1.3450 3.5950 1.6150 ;
      END
   END C
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 2.2950 0.1050 2.6250 0.5800 ;
	    RECT 3.2150 0.1050 3.5950 1.1050 ;
	    RECT 2.2950 0.0850 3.5950 0.1050 ;
	    RECT 0.0000 -0.0850 3.6800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.6800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.6800 3.4850 ;
	    RECT 0.0900 3.2950 3.5950 3.3150 ;
	    RECT 0.0900 1.8700 0.3450 3.2950 ;
	    RECT 1.0150 2.2950 1.1850 3.2950 ;
	    RECT 1.8550 2.2950 2.5450 3.2950 ;
	    RECT 3.2150 1.8050 3.5950 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.6800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0900 0.5800 0.3450 0.9350 ;
	    RECT 1.3550 0.7950 3.0450 1.1300 ;
	    RECT 0.0900 0.3700 2.1050 0.5800 ;
   END
END efs8hd_nand3_2
MACRO efs8hd_nand3b_2
   CLASS CORE ;
   FOREIGN efs8hd_nand3b_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.1400 BY 3.4000 ;
   SITE unitehd ;
   PIN AN
      PORT
         LAYER li1 ;
	    RECT 0.4300 1.3450 0.7800 1.6150 ;
      END
   END AN
   PIN C
      PORT
         LAYER li1 ;
	    RECT 1.0600 1.3450 1.7400 1.6150 ;
      END
   END C
   PIN B
      PORT
         LAYER li1 ;
	    RECT 1.9500 1.3450 3.1400 1.6150 ;
      END
   END B
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 1.0600 2.5050 1.3900 3.0800 ;
	    RECT 1.9000 2.5050 2.2300 3.0800 ;
	    RECT 1.0600 2.4450 2.2300 2.5050 ;
	    RECT 3.2600 2.5050 3.5100 3.0800 ;
	    RECT 3.2600 2.4450 4.0500 2.5050 ;
	    RECT 1.0600 2.2300 4.0500 2.4450 ;
	    RECT 3.8500 1.1300 4.0500 2.2300 ;
	    RECT 3.2600 0.7950 4.0500 1.1300 ;
      END
   END Y
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5800 0.1050 0.8900 1.1300 ;
	    RECT 1.5600 0.1050 1.8100 0.6800 ;
	    RECT 0.5800 0.0850 1.8100 0.1050 ;
	    RECT 0.0000 -0.0850 4.1400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.1400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.1400 3.4850 ;
	    RECT 0.5800 3.2950 4.0500 3.3150 ;
	    RECT 0.5800 2.2950 0.8900 3.2950 ;
	    RECT 1.5600 2.7200 1.7300 3.2950 ;
	    RECT 2.4000 2.7200 2.6500 3.2950 ;
	    RECT 2.8400 2.7200 3.0900 3.2950 ;
	    RECT 3.7600 2.7200 4.0500 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.1400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0900 2.5800 0.4100 3.0800 ;
	    RECT 0.0900 2.0200 0.2600 2.5800 ;
	    RECT 0.0900 1.8050 3.6500 2.0200 ;
	    RECT 0.0900 0.8200 0.2600 1.8050 ;
	    RECT 3.3200 1.3450 3.6500 1.8050 ;
	    RECT 1.0600 0.8950 2.7500 1.1300 ;
	    RECT 0.0900 0.3200 0.4100 0.8200 ;
	    RECT 1.0600 0.3200 1.3900 0.8950 ;
	    RECT 2.0000 0.7950 2.7500 0.8950 ;
	    RECT 2.9200 0.5800 3.0900 1.1300 ;
	    RECT 2.0000 0.3200 4.0500 0.5800 ;
   END
END efs8hd_nand3b_2
MACRO efs8hd_o2111ai_2
   CLASS CORE ;
   FOREIGN efs8hd_o2111ai_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.5200 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.6050 2.0800 0.8650 3.0800 ;
	    RECT 1.5350 2.0800 1.7250 3.0800 ;
	    RECT 2.3950 2.0800 2.5750 3.0800 ;
	    RECT 3.8150 2.0800 4.0050 2.6300 ;
	    RECT 0.6050 1.8700 4.0050 2.0800 ;
	    RECT 0.6050 1.1300 0.8650 1.8700 ;
	    RECT 0.6050 0.7700 0.9350 1.1300 ;
      END
   END Y
   PIN D1
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3450 0.4250 1.6950 ;
      END
   END D1
   PIN C1
      PORT
         LAYER li1 ;
	    RECT 1.0450 1.3450 1.7900 1.6550 ;
      END
   END C1
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 2.2000 1.3450 3.1850 1.6550 ;
      END
   END B1
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 3.3650 1.3450 4.4550 1.6550 ;
      END
   END A2
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 4.6350 1.3450 5.4350 1.6550 ;
      END
   END A1
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 3.7400 0.1050 4.0700 0.6050 ;
	    RECT 4.6000 0.1050 4.9300 0.6000 ;
	    RECT 3.7400 0.0850 4.9300 0.1050 ;
	    RECT 0.0000 -0.0850 5.5200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.5200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.5200 3.4850 ;
	    RECT 0.1750 3.2950 4.9300 3.3150 ;
	    RECT 0.1750 1.9050 0.4250 3.2950 ;
	    RECT 1.0350 2.2950 1.3650 3.2950 ;
	    RECT 1.8950 2.3000 2.2250 3.2950 ;
	    RECT 2.7550 2.2950 3.0850 3.2950 ;
	    RECT 4.6700 2.3200 4.9300 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.5200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 3.3100 2.8450 4.5000 3.0800 ;
	    RECT 3.3100 2.2950 3.5700 2.8450 ;
	    RECT 4.2400 2.1050 4.5000 2.8450 ;
	    RECT 5.1000 2.1050 5.3600 3.0800 ;
	    RECT 4.2400 1.8950 5.3600 2.1050 ;
	    RECT 0.1750 0.5550 0.4350 1.0800 ;
	    RECT 1.1150 0.9200 2.2750 1.1300 ;
	    RECT 1.1150 0.5550 1.3000 0.9200 ;
	    RECT 1.9250 0.7750 2.2750 0.9200 ;
	    RECT 2.4500 0.8200 5.4350 1.0500 ;
	    RECT 0.1750 0.3250 1.3000 0.5550 ;
	    RECT 1.4700 0.6650 1.7600 0.7050 ;
	    RECT 1.4700 0.5550 1.7750 0.6650 ;
	    RECT 2.8800 0.5550 3.2100 0.6050 ;
	    RECT 1.4700 0.3200 3.2100 0.5550 ;
	    RECT 3.3800 0.4550 3.5700 0.8200 ;
	    RECT 4.2400 0.8150 5.4350 0.8200 ;
	    RECT 4.2400 0.4550 4.4300 0.8150 ;
	    RECT 5.1000 0.4550 5.4350 0.8150 ;
   END
END efs8hd_o2111ai_2
MACRO efs8hd_o211ai_2
   CLASS CORE ;
   FOREIGN efs8hd_o211ai_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.6000 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5450 2.1400 0.8050 3.0800 ;
	    RECT 1.4750 2.1400 1.6650 3.0800 ;
	    RECT 2.8250 2.1400 3.1550 2.6550 ;
	    RECT 0.5450 1.9250 3.1550 2.1400 ;
	    RECT 0.5450 0.8400 0.8750 1.9250 ;
      END
   END Y
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 3.7050 1.2900 4.4550 1.6200 ;
	    RECT 4.1150 0.9550 4.4550 1.2900 ;
      END
   END A1
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 1.0450 1.3450 1.9050 1.7050 ;
      END
   END B1
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 2.3650 1.3450 3.5350 1.6950 ;
      END
   END A2
   PIN C1
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.2450 0.3750 2.4650 ;
      END
   END C1
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 2.3950 0.1050 2.7250 0.5550 ;
	    RECT 3.2550 0.1050 3.5850 0.5550 ;
	    RECT 4.1150 0.1050 4.4450 0.5550 ;
	    RECT 2.3950 0.0850 4.4450 0.1050 ;
	    RECT 0.0000 -0.0850 4.6000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.6000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.6000 3.4850 ;
	    RECT 0.1150 3.2950 4.0150 3.3150 ;
	    RECT 0.1150 2.7200 0.3750 3.2950 ;
	    RECT 0.9750 2.3950 1.3050 3.2950 ;
	    RECT 1.8350 2.3950 2.1650 3.2950 ;
	    RECT 3.6850 2.3300 4.0150 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.6000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 2.3950 2.8700 3.5150 3.0800 ;
	    RECT 2.3950 2.6250 2.6550 2.8700 ;
	    RECT 3.3250 2.1200 3.5150 2.8700 ;
	    RECT 4.1850 2.1200 4.4450 3.0800 ;
	    RECT 3.3250 1.9050 4.4450 2.1200 ;
	    RECT 1.0450 0.5800 1.2350 1.1150 ;
	    RECT 1.4050 0.7950 3.9450 1.0550 ;
	    RECT 3.7550 0.6450 3.9450 0.7950 ;
	    RECT 1.0450 0.5550 2.1650 0.5800 ;
	    RECT 0.0950 0.3200 2.1650 0.5550 ;
   END
END efs8hd_o211ai_2
MACRO efs8hd_o21ai_2
   CLASS CORE ;
   FOREIGN efs8hd_o21ai_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.2200 BY 3.4000 ;
   SITE unitehd ;
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 2.8150 0.7650 3.1300 1.7500 ;
      END
   END B1
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 0.1200 1.7850 2.0950 2.0200 ;
	    RECT 0.1200 1.3050 0.4350 1.7850 ;
	    RECT 1.6000 1.3450 2.0950 1.7850 ;
      END
   END A1
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 0.6050 1.3450 1.4200 1.6150 ;
      END
   END A2
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.9950 2.4550 1.2950 2.6550 ;
	    RECT 2.4100 2.4550 2.6450 3.0800 ;
	    RECT 0.9950 2.2300 2.6450 2.4550 ;
	    RECT 2.4350 0.7450 2.6450 2.2300 ;
      END
   END Y
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.6150 0.1050 0.7850 0.6800 ;
	    RECT 1.5250 0.1050 1.6950 0.6800 ;
	    RECT 0.6150 0.0850 1.6950 0.1050 ;
	    RECT 0.0000 -0.0850 3.2200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.2200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.2200 3.4850 ;
	    RECT 0.1050 3.2950 3.1250 3.3150 ;
	    RECT 0.1050 2.2300 0.4350 3.2950 ;
	    RECT 1.9100 2.7200 2.2400 3.2950 ;
	    RECT 2.8150 1.9650 3.1250 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.2200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.6050 2.8700 1.7150 3.0800 ;
	    RECT 0.6050 2.2300 0.8250 2.8700 ;
	    RECT 1.5250 2.6700 1.7150 2.8700 ;
	    RECT 0.1050 0.8950 2.2650 1.1050 ;
	    RECT 0.1050 0.3200 0.4350 0.8950 ;
	    RECT 0.9650 0.3200 1.2950 0.8950 ;
	    RECT 1.9350 0.5300 2.2650 0.8950 ;
	    RECT 2.7950 0.5300 3.1250 0.5950 ;
	    RECT 1.9350 0.3200 3.1250 0.5300 ;
   END
END efs8hd_o21ai_2
MACRO efs8hd_o21bai_2
   CLASS CORE ;
   FOREIGN efs8hd_o21bai_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.1400 BY 3.4000 ;
   SITE unitehd ;
   PIN B1N
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.1050 0.4950 1.6550 ;
      END
   END B1N
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 1.9500 1.3450 3.0900 1.6150 ;
      END
   END A2
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 3.2600 1.3450 4.0550 1.6150 ;
      END
   END A1
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 1.0850 2.0200 1.2550 3.0800 ;
	    RECT 2.4050 2.0200 2.6500 2.6550 ;
	    RECT 1.0850 1.8050 2.6500 2.0200 ;
	    RECT 1.5250 1.1300 1.7800 1.8050 ;
	    RECT 1.5250 0.8050 1.8550 1.1300 ;
      END
   END Y
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1800 0.1050 0.3500 0.9350 ;
	    RECT 2.4450 0.1050 2.6150 0.6950 ;
	    RECT 3.2850 0.1050 3.4550 0.6950 ;
	    RECT 0.1800 0.0850 3.4550 0.1050 ;
	    RECT 0.0000 -0.0850 4.1400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.1400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.1400 3.4850 ;
	    RECT 0.5850 3.2950 3.5350 3.3150 ;
	    RECT 0.5850 2.3450 0.9150 3.2950 ;
	    RECT 1.4700 2.2450 1.7200 3.2950 ;
	    RECT 3.2050 2.2950 3.5350 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.1400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 1.9550 2.8700 3.0350 3.0800 ;
	    RECT 0.1800 2.0800 0.3500 2.3950 ;
	    RECT 1.9550 2.2450 2.2350 2.8700 ;
	    RECT 2.8650 2.0800 3.0350 2.8700 ;
	    RECT 3.7050 2.0800 3.9800 3.0800 ;
	    RECT 0.1800 1.8700 0.8650 2.0800 ;
	    RECT 0.6950 1.5550 0.8650 1.8700 ;
	    RECT 2.8650 1.8200 3.9800 2.0800 ;
	    RECT 0.6950 1.3450 1.3350 1.5550 ;
	    RECT 0.6950 0.9700 0.8650 1.3450 ;
	    RECT 0.6000 0.5550 0.8650 0.9700 ;
	    RECT 1.0750 0.5950 1.3550 1.1300 ;
	    RECT 2.0250 0.9050 3.9800 1.1300 ;
	    RECT 2.0250 0.5950 2.2750 0.9050 ;
	    RECT 1.0750 0.3200 2.2750 0.5950 ;
	    RECT 2.7850 0.3200 3.1150 0.9050 ;
	    RECT 3.6250 0.3300 3.9800 0.9050 ;
   END
END efs8hd_o21bai_2
MACRO efs8hd_o221ai_2
   CLASS CORE ;
   FOREIGN efs8hd_o221ai_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.5200 BY 3.4000 ;
   SITE unitehd ;
   PIN C1
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3450 0.4350 1.6150 ;
      END
   END C1
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 1.0200 1.8050 3.2600 2.0200 ;
	    RECT 1.0200 1.3450 2.0350 1.8050 ;
	    RECT 2.9250 1.3450 3.2600 1.8050 ;
      END
   END B1
   PIN B2
      PORT
         LAYER li1 ;
	    RECT 2.2050 1.3450 2.7550 1.6150 ;
      END
   END B2
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 3.8250 1.3450 4.4750 1.6150 ;
      END
   END A2
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 3.4300 1.7850 4.8150 2.0200 ;
	    RECT 3.4300 1.3050 3.6550 1.7850 ;
	    RECT 4.6450 1.6150 4.8150 1.7850 ;
	    RECT 4.6450 1.3450 5.4350 1.6150 ;
      END
   END A1
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5600 2.4450 0.8100 3.0800 ;
	    RECT 2.3400 2.4450 2.5900 2.6550 ;
	    RECT 4.1000 2.4450 4.3500 2.6550 ;
	    RECT 0.5600 2.2300 4.3500 2.4450 ;
	    RECT 0.5600 1.8050 0.8450 2.2300 ;
	    RECT 0.6050 1.0800 0.8450 1.8050 ;
	    RECT 0.5150 0.8050 0.8450 1.0800 ;
      END
   END Y
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 3.7200 0.1050 3.8900 0.6950 ;
	    RECT 4.5600 0.1050 4.7300 0.6950 ;
	    RECT 3.7200 0.0850 4.7300 0.1050 ;
	    RECT 0.0000 -0.0850 5.5200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.5200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.5200 3.4850 ;
	    RECT 0.1400 3.2950 5.1900 3.3150 ;
	    RECT 0.1400 1.8200 0.3900 3.2950 ;
	    RECT 0.9800 2.6550 1.7500 3.2950 ;
	    RECT 3.1800 2.6550 3.5100 3.2950 ;
	    RECT 4.9850 1.8200 5.1900 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.5200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 1.9200 2.8700 3.0100 3.0800 ;
	    RECT 1.9200 2.6550 2.1700 2.8700 ;
	    RECT 2.7600 2.6550 3.0100 2.8700 ;
	    RECT 3.6800 2.8700 4.7700 3.0800 ;
	    RECT 3.6800 2.6550 3.9300 2.8700 ;
	    RECT 4.5200 2.2300 4.7700 2.8700 ;
	    RECT 0.1000 0.5950 0.3450 1.1200 ;
	    RECT 1.0150 0.8050 3.0500 1.1300 ;
	    RECT 3.2200 0.9200 5.2300 1.1300 ;
	    RECT 1.0150 0.5950 1.2700 0.8050 ;
	    RECT 3.2200 0.5950 3.5500 0.9200 ;
	    RECT 0.1000 0.3200 1.2700 0.5950 ;
	    RECT 1.4550 0.3200 3.5500 0.5950 ;
	    RECT 4.0600 0.9050 5.2300 0.9200 ;
	    RECT 4.0600 0.3200 4.3900 0.9050 ;
	    RECT 4.9000 0.3200 5.2300 0.9050 ;
   END
END efs8hd_o221ai_2
MACRO efs8hd_o22ai_2
   CLASS CORE ;
   FOREIGN efs8hd_o22ai_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.6000 BY 3.4000 ;
   SITE unitehd ;
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 0.1450 1.3000 0.8950 1.6300 ;
      END
   END B1
   PIN B2
      PORT
         LAYER li1 ;
	    RECT 1.0650 1.3450 1.9250 1.6150 ;
      END
   END B2
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 2.4450 1.3050 3.1950 1.6350 ;
      END
   END A2
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 3.3650 1.3450 4.1650 1.6150 ;
      END
   END A1
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 1.4150 2.0300 1.6650 2.6550 ;
	    RECT 2.8150 2.0300 3.0750 2.6550 ;
	    RECT 1.4150 1.8050 3.0750 2.0300 ;
	    RECT 1.4150 1.7850 2.2750 1.8050 ;
	    RECT 2.0950 1.1300 2.2750 1.7850 ;
	    RECT 0.5350 0.9050 2.2750 1.1300 ;
	    RECT 0.5350 0.8050 0.8650 0.9050 ;
	    RECT 1.3750 0.8050 1.7050 0.9050 ;
      END
   END Y
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 2.8550 0.1050 3.0250 0.6950 ;
	    RECT 3.6950 0.1050 3.8650 0.6950 ;
	    RECT 2.8550 0.0850 3.8650 0.1050 ;
	    RECT 0.0000 -0.0850 4.6000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.6000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.6000 3.4850 ;
	    RECT 0.5750 3.2950 3.9050 3.3150 ;
	    RECT 0.5750 2.2450 0.8250 3.2950 ;
	    RECT 3.6550 2.2450 3.9050 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.6000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1500 2.0300 0.4050 3.0800 ;
	    RECT 0.9950 2.8700 2.0850 3.0800 ;
	    RECT 0.9950 2.0300 1.2450 2.8700 ;
	    RECT 1.8350 2.2450 2.0850 2.8700 ;
	    RECT 2.3950 2.8700 3.4850 3.0800 ;
	    RECT 2.3950 2.2450 2.6450 2.8700 ;
	    RECT 0.1500 1.8200 1.2450 2.0300 ;
	    RECT 3.2450 2.0300 3.4850 2.8700 ;
	    RECT 4.0750 2.0300 4.3300 3.0800 ;
	    RECT 3.2450 1.8200 4.3300 2.0300 ;
	    RECT 0.0900 0.5950 0.3650 1.1300 ;
	    RECT 2.5100 0.9050 4.3650 1.1300 ;
	    RECT 2.5100 0.5950 2.6800 0.9050 ;
	    RECT 0.0900 0.3800 2.6800 0.5950 ;
	    RECT 3.1950 0.3200 3.5250 0.9050 ;
	    RECT 4.0350 0.3200 4.3650 0.9050 ;
   END
END efs8hd_o22ai_2
MACRO efs8hd_o2bb2ai_2
   CLASS CORE ;
   FOREIGN efs8hd_o2bb2ai_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.5200 BY 3.4000 ;
   SITE unitehd ;
   PIN A1N
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.7850 1.9450 2.0200 ;
	    RECT 0.0900 1.3050 0.4350 1.7850 ;
	    RECT 1.6150 1.3450 1.9450 1.7850 ;
      END
   END A1N
   PIN A2N
      PORT
         LAYER li1 ;
	    RECT 0.6050 1.3450 1.4000 1.6150 ;
      END
   END A2N
   PIN B2
      PORT
         LAYER li1 ;
	    RECT 3.8250 1.3450 4.5000 1.6150 ;
      END
   END B2
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 3.4100 1.8050 5.4350 2.0200 ;
	    RECT 3.4100 1.3050 3.6550 1.8050 ;
	    RECT 4.7300 1.3450 5.4350 1.8050 ;
      END
   END B1
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 2.7450 2.4450 3.0350 3.0800 ;
	    RECT 4.0800 2.4450 4.3300 2.6550 ;
	    RECT 2.7450 2.2300 4.3300 2.4450 ;
	    RECT 2.7450 1.3450 3.2150 2.2300 ;
	    RECT 2.7450 0.8050 3.0750 1.3450 ;
      END
   END Y
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1950 0.1050 0.3650 1.1200 ;
	    RECT 1.8750 0.1050 2.0450 0.6950 ;
	    RECT 3.7000 0.1050 3.8700 0.6950 ;
	    RECT 4.5400 0.1050 4.7100 0.6950 ;
	    RECT 0.1950 0.0850 4.7100 0.1050 ;
	    RECT 0.0000 -0.0850 5.5200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.5200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.5200 3.4850 ;
	    RECT 0.1500 3.2950 5.1700 3.3150 ;
	    RECT 0.1500 2.2450 0.4000 3.2950 ;
	    RECT 0.9950 2.6700 1.2450 3.2950 ;
	    RECT 1.8350 2.6700 2.5750 3.2950 ;
	    RECT 3.2050 2.6550 3.4900 3.2950 ;
	    RECT 4.9650 2.2450 5.1700 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.5200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.5750 2.4550 0.8250 3.0800 ;
	    RECT 3.6600 2.8700 4.7500 3.0800 ;
	    RECT 3.6600 2.6550 3.9100 2.8700 ;
	    RECT 1.4150 2.4550 1.6650 2.6550 ;
	    RECT 0.5750 2.2300 2.2850 2.4550 ;
	    RECT 4.5000 2.2300 4.7500 2.8700 ;
	    RECT 2.1150 1.6550 2.2850 2.2300 ;
	    RECT 2.1150 1.2450 2.5750 1.6550 ;
	    RECT 2.1150 1.1300 2.2850 1.2450 ;
	    RECT 0.5350 0.5950 0.7850 1.1200 ;
	    RECT 0.9550 0.9050 2.2850 1.1300 ;
	    RECT 3.2450 0.9200 5.2100 1.1300 ;
	    RECT 0.9550 0.8050 1.2850 0.9050 ;
	    RECT 2.3250 0.5950 2.5750 0.6950 ;
	    RECT 3.2450 0.5950 3.5300 0.9200 ;
	    RECT 0.5350 0.3800 1.7050 0.5950 ;
	    RECT 2.3250 0.3200 3.5300 0.5950 ;
	    RECT 4.0400 0.9050 5.2100 0.9200 ;
	    RECT 4.0400 0.3200 4.3700 0.9050 ;
	    RECT 4.8800 0.3200 5.2100 0.9050 ;
   END
END efs8hd_o2bb2ai_2
MACRO efs8hd_o311ai_2
   CLASS CORE ;
   FOREIGN efs8hd_o311ai_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.9800 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 2.4150 2.1550 2.6650 2.6550 ;
	    RECT 3.3350 2.1550 3.5050 3.0800 ;
	    RECT 4.5150 2.1550 4.8250 3.0800 ;
	    RECT 5.4950 2.1550 5.8950 3.0800 ;
	    RECT 2.4150 1.8550 5.8950 2.1550 ;
	    RECT 4.6250 1.1050 4.9150 1.8550 ;
	    RECT 4.6250 0.8050 5.8950 1.1050 ;
	    RECT 5.5150 0.3200 5.8950 0.8050 ;
      END
   END Y
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3200 1.2350 1.6450 ;
      END
   END A1
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 1.4050 1.3050 2.1550 1.6450 ;
      END
   END A2
   PIN A3
      PORT
         LAYER li1 ;
	    RECT 2.3250 1.3200 3.0750 1.6450 ;
      END
   END A3
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 3.3650 1.3200 4.4550 1.6450 ;
      END
   END B1
   PIN C1
      PORT
         LAYER li1 ;
	    RECT 5.0850 1.3200 5.8950 1.6450 ;
      END
   END C1
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.6550 0.1050 0.9850 0.6050 ;
	    RECT 1.4950 0.1050 1.8250 0.6050 ;
	    RECT 2.3350 0.1050 3.1050 0.6050 ;
	    RECT 0.6550 0.0850 3.1050 0.1050 ;
	    RECT 0.0000 -0.0850 5.9800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.9800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.9800 3.4850 ;
	    RECT 0.6350 3.2950 5.3250 3.3150 ;
	    RECT 0.6350 2.3700 0.9650 3.2950 ;
	    RECT 3.6750 2.3700 4.3450 3.2950 ;
	    RECT 4.9950 2.3700 5.3250 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.9800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.1550 0.4650 3.0800 ;
	    RECT 1.1350 2.1550 1.3050 3.0800 ;
	    RECT 1.4750 2.8700 3.1650 3.0800 ;
	    RECT 1.4750 2.3700 1.8050 2.8700 ;
	    RECT 1.9750 2.1550 2.2250 2.6550 ;
	    RECT 2.8350 2.3700 3.1650 2.8700 ;
	    RECT 0.0850 1.8550 2.2250 2.1550 ;
	    RECT 0.0850 0.8200 4.3850 1.1050 ;
	    RECT 0.0850 0.3200 0.4850 0.8200 ;
	    RECT 1.1550 0.3200 1.3250 0.8200 ;
	    RECT 1.9950 0.3200 2.1650 0.8200 ;
	    RECT 3.2750 0.3200 3.4450 0.8200 ;
	    RECT 3.6150 0.3200 5.3450 0.6050 ;
   END
END efs8hd_o311ai_2
MACRO efs8hd_o31ai_2
   CLASS CORE ;
   FOREIGN efs8hd_o31ai_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.6000 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 2.3350 2.0800 2.6650 2.6550 ;
	    RECT 3.1750 2.0800 3.5050 3.0800 ;
	    RECT 4.1750 2.0800 4.5150 3.0800 ;
	    RECT 2.3350 1.8700 4.5150 2.0800 ;
	    RECT 3.6750 0.7450 4.0050 1.8700 ;
      END
   END Y
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 4.1750 0.7650 4.5150 1.6550 ;
      END
   END B1
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.3200 1.2400 1.6550 ;
      END
   END A1
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 1.4100 1.3200 2.2200 1.6550 ;
      END
   END A2
   PIN A3
      PORT
         LAYER li1 ;
	    RECT 2.3900 1.3200 3.2050 1.6550 ;
      END
   END A3
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.6150 0.1050 0.7850 0.6800 ;
	    RECT 1.4550 0.1050 1.9650 0.6800 ;
	    RECT 2.6750 0.1050 3.0050 0.6800 ;
	    RECT 0.6150 0.0850 3.0050 0.1050 ;
	    RECT 0.0000 -0.0850 4.6000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.6000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.6000 3.4850 ;
	    RECT 0.6150 3.2950 4.0050 3.3150 ;
	    RECT 0.6150 2.2950 0.7850 3.2950 ;
	    RECT 3.6750 2.2950 4.0050 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.6000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0900 2.0800 0.4450 3.0800 ;
	    RECT 0.9550 2.0800 1.2850 3.0800 ;
	    RECT 1.4550 2.8700 3.0050 3.0800 ;
	    RECT 1.4550 2.2950 1.6250 2.8700 ;
	    RECT 1.7950 2.0800 2.1250 2.6550 ;
	    RECT 2.8350 2.2950 3.0050 2.8700 ;
	    RECT 0.0900 1.8700 2.1250 2.0800 ;
	    RECT 0.0900 0.8950 3.5050 1.1050 ;
	    RECT 0.0900 0.3200 0.4450 0.8950 ;
	    RECT 0.9550 0.3200 1.2850 0.8950 ;
	    RECT 2.1750 0.3200 2.5050 0.8950 ;
	    RECT 3.1750 0.5300 3.5050 0.8950 ;
	    RECT 4.1350 0.5300 4.5150 0.5950 ;
	    RECT 3.1750 0.3200 4.5150 0.5300 ;
   END
END efs8hd_o31ai_2
MACRO efs8hd_o32ai_2
   CLASS CORE ;
   FOREIGN efs8hd_o32ai_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.9800 BY 3.4000 ;
   SITE unitehd ;
   PIN B2
      PORT
         LAYER li1 ;
	    RECT 0.0900 1.3450 0.8450 1.6550 ;
      END
   END B2
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 1.0150 1.3450 1.7050 1.6550 ;
      END
   END B1
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5150 2.0800 0.8450 2.6200 ;
	    RECT 2.7750 2.0800 3.1050 2.6050 ;
	    RECT 0.5150 1.8700 3.1050 2.0800 ;
	    RECT 1.8750 1.3800 2.1700 1.8700 ;
	    RECT 1.8750 1.1300 2.0450 1.3800 ;
	    RECT 0.5150 0.8200 2.0450 1.1300 ;
      END
   END Y
   PIN A3
      PORT
         LAYER li1 ;
	    RECT 2.4050 1.3450 3.0750 1.6550 ;
      END
   END A3
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 3.3650 1.3450 4.4800 1.6550 ;
      END
   END A2
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 4.7450 1.3450 5.8650 1.6550 ;
      END
   END A1
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 2.6200 0.1050 2.9500 0.6800 ;
	    RECT 3.6350 0.1050 3.8050 0.6800 ;
	    RECT 4.9050 0.1050 5.2350 0.6800 ;
	    RECT 2.6200 0.0850 5.2350 0.1050 ;
	    RECT 0.0000 -0.0850 5.9800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.9800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.9800 3.4850 ;
	    RECT 1.4350 3.2950 5.7150 3.3150 ;
	    RECT 1.4350 2.7200 1.6050 3.2950 ;
	    RECT 4.6200 2.2950 4.8250 3.2950 ;
	    RECT 5.4950 1.8700 5.7150 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.9800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0900 2.8700 1.2650 3.0800 ;
	    RECT 0.0900 1.8700 0.3450 2.8700 ;
	    RECT 1.0150 2.5050 1.2650 2.8700 ;
	    RECT 1.7750 2.5050 2.1050 3.0700 ;
	    RECT 1.0150 2.2950 2.1050 2.5050 ;
	    RECT 2.3350 2.8200 4.3850 3.0550 ;
	    RECT 2.3350 2.2950 2.5850 2.8200 ;
	    RECT 3.2750 1.8700 3.4450 2.8200 ;
	    RECT 3.6150 2.0800 3.9450 2.6050 ;
	    RECT 4.1350 2.2950 4.3850 2.8200 ;
	    RECT 4.9950 2.0800 5.3250 3.0750 ;
	    RECT 3.6150 1.8700 5.3250 2.0800 ;
	    RECT 0.0900 0.6050 0.3450 1.1300 ;
	    RECT 2.2350 0.8950 5.7550 1.1300 ;
	    RECT 2.2350 0.6050 2.4050 0.8950 ;
	    RECT 0.0900 0.3200 2.4050 0.6050 ;
	    RECT 3.1350 0.3200 3.4650 0.8950 ;
	    RECT 4.0550 0.3200 4.7250 0.8950 ;
	    RECT 5.4250 0.3200 5.7550 0.8950 ;
   END
END efs8hd_o32ai_2
MACRO efs8hd_o41ai_2
   CLASS CORE ;
   FOREIGN efs8hd_o41ai_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.9800 BY 3.4000 ;
   SITE unitehd ;
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 0.5150 2.0800 0.8450 3.0800 ;
	    RECT 1.8750 2.0800 2.2050 2.6550 ;
	    RECT 0.5150 1.8800 2.2050 2.0800 ;
	    RECT 0.6100 1.8050 2.2050 1.8800 ;
	    RECT 0.6100 1.1050 0.8450 1.8050 ;
	    RECT 0.5150 0.7950 0.8450 1.1050 ;
      END
   END Y
   PIN B1
      PORT
         LAYER li1 ;
	    RECT 0.1050 1.3450 0.4400 1.6150 ;
      END
   END B1
   PIN A4
      PORT
         LAYER li1 ;
	    RECT 1.5000 1.3050 2.2750 1.6350 ;
      END
   END A4
   PIN A3
      PORT
         LAYER li1 ;
	    RECT 2.4450 1.3450 3.5800 1.6150 ;
      END
   END A3
   PIN A2
      PORT
         LAYER li1 ;
	    RECT 3.7800 1.3450 4.5400 1.6150 ;
      END
   END A2
   PIN A1
      PORT
         LAYER li1 ;
	    RECT 4.7200 1.3450 5.8950 1.6150 ;
      END
   END A1
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 1.4550 0.1050 1.7050 0.6800 ;
	    RECT 2.3750 0.1050 2.5450 0.6800 ;
	    RECT 3.2150 0.1050 3.4500 0.6800 ;
	    RECT 4.1950 0.1050 4.3650 0.6800 ;
	    RECT 5.0350 0.1050 5.2050 0.6800 ;
	    RECT 1.4550 0.0850 5.2050 0.1050 ;
	    RECT 0.0000 -0.0850 5.9800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.9800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.9800 3.4850 ;
	    RECT 0.0850 3.2950 5.2850 3.3150 ;
	    RECT 0.0850 1.8700 0.3450 3.2950 ;
	    RECT 1.0150 2.2950 1.2650 3.2950 ;
	    RECT 4.9550 2.2300 5.2850 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.9800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 1.4550 2.8700 2.5450 3.0800 ;
	    RECT 1.4550 2.2950 1.7050 2.8700 ;
	    RECT 2.3750 2.0200 2.5450 2.8700 ;
	    RECT 2.7150 2.8700 4.4450 3.0800 ;
	    RECT 2.7150 2.2950 3.0450 2.8700 ;
	    RECT 3.2150 2.0200 3.4650 2.6550 ;
	    RECT 2.3750 1.8050 3.4650 2.0200 ;
	    RECT 3.6950 2.0200 3.9450 2.6550 ;
	    RECT 4.1150 2.2950 4.4450 2.8700 ;
	    RECT 4.6150 2.0200 4.7850 3.0800 ;
	    RECT 5.4550 2.0200 5.7050 3.0800 ;
	    RECT 3.6950 1.8050 5.7050 2.0200 ;
	    RECT 0.0850 0.5800 0.3450 1.1300 ;
	    RECT 1.0150 0.9200 5.7050 1.1300 ;
	    RECT 1.0150 0.5800 1.2650 0.9200 ;
	    RECT 0.0850 0.3200 1.2650 0.5800 ;
	    RECT 1.8750 0.3200 2.2050 0.9200 ;
	    RECT 2.7150 0.3200 3.0450 0.9200 ;
	    RECT 3.6950 0.3200 4.0250 0.9200 ;
	    RECT 4.5350 0.3200 4.8650 0.9200 ;
	    RECT 5.3750 0.3200 5.7050 0.9200 ;
   END
END efs8hd_o41ai_2
MACRO efs8hd_or2_2
   CLASS CORE ;
   FOREIGN efs8hd_or2_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 2.3000 BY 3.4000 ;
   SITE unitehd ;
   PIN B
      PORT
         LAYER li1 ;
	    RECT 0.1450 0.7650 0.3450 1.6550 ;
      END
   END B
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.8650 0.7650 1.2750 1.6550 ;
      END
   END A
   PIN X
      PORT
         LAYER li1 ;
	    RECT 1.4400 2.5050 1.7700 3.0800 ;
	    RECT 1.4400 2.2950 2.2150 2.5050 ;
	    RECT 1.7850 1.0300 2.2150 2.2950 ;
	    RECT 1.5200 0.8200 2.2150 1.0300 ;
	    RECT 1.5200 0.4800 1.6900 0.8200 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1050 0.1050 0.3450 0.5950 ;
	    RECT 1.0150 0.1050 1.3500 0.5950 ;
	    RECT 1.8600 0.1050 2.1900 0.6050 ;
	    RECT 0.1050 0.0850 2.1900 0.1050 ;
	    RECT 0.0000 -0.0850 2.3000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 2.3000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 2.3000 3.4850 ;
	    RECT 1.1000 3.2950 2.1100 3.3150 ;
	    RECT 1.1000 2.2950 1.2700 3.2950 ;
	    RECT 1.9400 2.7200 2.1100 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 2.3000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1550 2.0800 0.5150 2.3000 ;
	    RECT 0.1550 1.8700 1.6150 2.0800 ;
	    RECT 0.5150 0.5950 0.6950 1.8700 ;
	    RECT 1.4450 1.2450 1.6150 1.8700 ;
	    RECT 0.5150 0.3200 0.8450 0.5950 ;
   END
END efs8hd_or2_2
MACRO efs8hd_or2b_2
   CLASS CORE ;
   FOREIGN efs8hd_or2b_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.2200 BY 3.4000 ;
   SITE unitehd ;
   PIN BN
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3450 0.4250 1.6550 ;
      END
   END BN
   PIN X
      PORT
         LAYER li1 ;
	    RECT 2.4000 1.8700 2.6300 3.0800 ;
	    RECT 2.4600 0.9500 2.6300 1.8700 ;
	    RECT 2.4000 0.5200 2.6300 0.9500 ;
      END
   END X
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.5400 2.6050 1.7300 3.0200 ;
      END
   END A
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5900 0.1050 1.3200 0.7050 ;
	    RECT 1.8300 0.1050 2.2100 0.6050 ;
	    RECT 2.8000 0.1050 3.0550 1.1550 ;
	    RECT 0.5900 0.0850 3.0550 0.1050 ;
	    RECT 0.0000 -0.0850 3.2200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.2200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.2200 3.4850 ;
	    RECT 0.0850 3.2950 3.0550 3.3150 ;
	    RECT 0.0850 1.8700 0.3450 3.2950 ;
	    RECT 1.9100 2.2950 2.1900 3.2950 ;
	    RECT 2.8000 1.8250 3.0550 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.2200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.5950 1.6550 0.7650 2.3550 ;
	    RECT 0.9850 2.0800 1.4050 2.3950 ;
	    RECT 0.9850 1.8700 2.2300 2.0800 ;
	    RECT 2.0600 1.6550 2.2300 1.8700 ;
	    RECT 0.5950 1.2450 1.3300 1.6550 ;
	    RECT 2.0600 1.2450 2.2900 1.6550 ;
	    RECT 0.5950 1.1300 0.8400 1.2450 ;
	    RECT 0.1050 0.9200 0.8400 1.1300 ;
	    RECT 2.0600 1.0300 2.2300 1.2450 ;
	    RECT 0.1050 0.3300 0.4200 0.9200 ;
	    RECT 1.4900 0.8200 2.2300 1.0300 ;
	    RECT 1.4900 0.3800 1.6600 0.8200 ;
   END
END efs8hd_or2b_2
MACRO efs8hd_or3_2
   CLASS CORE ;
   FOREIGN efs8hd_or3_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 2.7600 BY 3.4000 ;
   SITE unitehd ;
   PIN C
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.1050 0.4350 1.6550 ;
      END
   END C
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.6050 1.6550 0.8300 2.0200 ;
	    RECT 0.6050 1.2450 1.4300 1.6550 ;
      END
   END A
   PIN X
      PORT
         LAYER li1 ;
	    RECT 1.9400 1.8700 2.2150 3.0800 ;
	    RECT 2.0450 0.9500 2.2150 1.8700 ;
	    RECT 1.9400 0.5200 2.2150 0.9500 ;
      END
   END X
   PIN B
      PORT
         LAYER li1 ;
	    RECT 0.0850 2.6550 1.2800 3.0200 ;
      END
   END B
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5300 0.1050 0.8600 0.5950 ;
	    RECT 1.3700 0.1050 1.7500 0.5950 ;
	    RECT 2.3850 0.1050 2.6750 1.1450 ;
	    RECT 0.5300 0.0850 2.6750 0.1050 ;
	    RECT 0.0000 -0.0850 2.7600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 2.7600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 2.7600 3.4850 ;
	    RECT 1.4500 3.2950 2.6750 3.3150 ;
	    RECT 1.4500 2.2950 1.7300 3.2950 ;
	    RECT 2.3850 1.7900 2.6750 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 2.7600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1050 2.2300 1.2700 2.4450 ;
	    RECT 0.1050 1.8700 0.4350 2.2300 ;
	    RECT 1.1000 2.0800 1.2700 2.2300 ;
	    RECT 1.1000 1.8700 1.7700 2.0800 ;
	    RECT 1.6000 1.6550 1.7700 1.8700 ;
	    RECT 1.6000 1.2450 1.8750 1.6550 ;
	    RECT 1.6000 0.9350 1.7700 1.2450 ;
	    RECT 0.1050 0.7650 1.7700 0.9350 ;
	    RECT 0.1050 0.3800 0.3600 0.7650 ;
	    RECT 1.0300 0.3800 1.2000 0.7650 ;
   END
END efs8hd_or3_2
MACRO efs8hd_or3b_2
   CLASS CORE ;
   FOREIGN efs8hd_or3b_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.2200 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 0.9350 1.7850 1.3300 2.2950 ;
	    RECT 0.9350 0.7450 1.1050 1.7850 ;
	    RECT 0.9350 0.3300 1.2850 0.7450 ;
      END
   END X
   PIN CN
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3450 0.4250 2.0500 ;
      END
   END CN
   PIN A
      PORT
         LAYER li1 ;
	    RECT 1.6950 1.3450 2.2300 2.0200 ;
      END
   END A
   PIN B
      PORT
         LAYER li1 ;
	    RECT 1.9350 2.6550 3.1350 2.9750 ;
      END
   END B
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5950 0.1050 0.7650 0.7050 ;
	    RECT 1.5200 0.1050 1.6900 0.7050 ;
	    RECT 2.3300 0.1050 2.6600 0.6050 ;
	    RECT 0.5950 0.0850 2.6600 0.1050 ;
	    RECT 0.0000 -0.0850 3.2200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.2200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.2200 3.4850 ;
	    RECT 0.5500 3.2950 1.7550 3.3150 ;
	    RECT 0.5500 2.8050 0.9100 3.2950 ;
	    RECT 1.4250 2.8050 1.7550 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.2200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.6350 0.3450 2.7750 ;
	    RECT 0.0850 2.4650 1.7200 2.6350 ;
	    RECT 0.0850 2.2650 0.7650 2.4650 ;
	    RECT 0.5950 1.1300 0.7650 2.2650 ;
	    RECT 1.5500 2.4450 1.7200 2.4650 ;
	    RECT 1.5500 2.2300 2.6600 2.4450 ;
	    RECT 2.4900 1.6550 2.6600 2.2300 ;
	    RECT 2.8300 1.8700 3.1350 2.4050 ;
	    RECT 0.0850 0.9200 0.7650 1.1300 ;
	    RECT 1.2750 1.1700 1.4450 1.6150 ;
	    RECT 2.4900 1.2450 2.7900 1.6550 ;
	    RECT 1.2750 1.1300 1.5950 1.1700 ;
	    RECT 1.2750 1.0300 2.1600 1.1300 ;
	    RECT 2.9650 1.0300 3.1350 1.8700 ;
	    RECT 1.2750 0.9550 3.1350 1.0300 ;
	    RECT 1.4250 0.9200 3.1350 0.9550 ;
	    RECT 0.0850 0.3650 0.3450 0.9200 ;
	    RECT 1.9900 0.8200 3.1350 0.9200 ;
	    RECT 1.9900 0.3800 2.1600 0.8200 ;
	    RECT 2.8300 0.7550 3.1350 0.8200 ;
	    RECT 2.8300 0.3800 3.0850 0.7550 ;
   END
END efs8hd_or3b_2
MACRO efs8hd_or4_2
   CLASS CORE ;
   FOREIGN efs8hd_or4_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.2200 BY 3.4000 ;
   SITE unitehd ;
   PIN D
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.7650 0.4350 1.6550 ;
      END
   END D
   PIN C
      PORT
         LAYER li1 ;
	    RECT 0.6050 1.2450 1.3200 2.0200 ;
      END
   END C
   PIN A
      PORT
         LAYER li1 ;
	    RECT 1.4900 1.1050 1.8950 1.6550 ;
      END
   END A
   PIN X
      PORT
         LAYER li1 ;
	    RECT 2.4050 1.8700 2.6800 3.0800 ;
	    RECT 2.5100 0.9500 2.6800 1.8700 ;
	    RECT 2.4050 0.5200 2.6800 0.9500 ;
      END
   END X
   PIN B
      PORT
         LAYER li1 ;
	    RECT 0.0850 2.6550 1.7450 3.0200 ;
      END
   END B
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0900 0.1050 0.4250 0.5950 ;
	    RECT 0.9950 0.1050 1.3250 0.5950 ;
	    RECT 1.8350 0.1050 2.2150 0.5950 ;
	    RECT 2.8500 0.1050 3.0200 1.2500 ;
	    RECT 0.0900 0.0850 3.0200 0.1050 ;
	    RECT 0.0000 -0.0850 3.2200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.2200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.2200 3.4850 ;
	    RECT 1.9150 3.2950 3.0200 3.3150 ;
	    RECT 1.9150 2.2950 2.1950 3.2950 ;
	    RECT 2.8500 1.8200 3.0200 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.2200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.2300 1.6800 2.4450 ;
	    RECT 0.0850 1.8700 0.4100 2.2300 ;
	    RECT 1.5100 2.0800 1.6800 2.2300 ;
	    RECT 1.5100 1.8700 2.2350 2.0800 ;
	    RECT 2.0650 1.6550 2.2350 1.8700 ;
	    RECT 2.0650 1.2450 2.3400 1.6550 ;
	    RECT 2.0650 0.9350 2.2350 1.2450 ;
	    RECT 0.6250 0.7650 2.2350 0.9350 ;
	    RECT 0.6250 0.3800 0.7950 0.7650 ;
	    RECT 1.4950 0.3800 1.6650 0.7650 ;
   END
END efs8hd_or4_2
MACRO efs8hd_or4b_2
   CLASS CORE ;
   FOREIGN efs8hd_or4b_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 3.6800 BY 3.4000 ;
   SITE unitehd ;
   PIN X
      PORT
         LAYER li1 ;
	    RECT 0.9350 1.8700 1.2500 2.2950 ;
	    RECT 0.9350 0.9900 1.1050 1.8700 ;
	    RECT 0.9350 0.8500 1.2450 0.9900 ;
	    RECT 0.9350 0.8450 1.2500 0.8500 ;
	    RECT 0.9700 0.3250 1.2500 0.8450 ;
      END
   END X
   PIN DN
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.3450 0.4250 1.9550 ;
      END
   END DN
   PIN A
      PORT
         LAYER li1 ;
	    RECT 1.7550 1.3450 2.2750 1.6150 ;
      END
   END A
   PIN C
      PORT
         LAYER li1 ;
	    RECT 2.4450 1.3450 3.5500 1.6150 ;
      END
   END C
   PIN B
      PORT
         LAYER li1 ;
	    RECT 1.9850 2.4650 2.6700 3.0200 ;
      END
   END B
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.6300 0.1050 0.8000 0.7050 ;
	    RECT 1.4350 0.1050 1.8150 0.6050 ;
	    RECT 2.3850 0.1050 2.7150 0.6050 ;
	    RECT 3.2250 0.1050 3.5550 0.7300 ;
	    RECT 0.6300 0.0850 3.5550 0.1050 ;
	    RECT 0.0000 -0.0850 3.6800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 3.6800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 3.6800 3.4850 ;
	    RECT 0.5150 3.2950 1.8150 3.3150 ;
	    RECT 0.5150 2.9200 0.8450 3.2950 ;
	    RECT 1.4800 2.9200 1.8150 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 3.6800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 2.8600 2.7700 3.3450 2.9800 ;
	    RECT 0.5100 2.4950 1.7150 2.7050 ;
	    RECT 0.5100 2.3650 0.7650 2.4950 ;
	    RECT 0.0850 2.1250 0.7650 2.3650 ;
	    RECT 1.4400 2.2950 1.7150 2.4950 ;
	    RECT 2.8600 2.2950 3.0300 2.7700 ;
	    RECT 1.4400 2.1250 3.0300 2.2950 ;
	    RECT 0.5950 1.1300 0.7650 2.1250 ;
	    RECT 3.2250 1.9550 3.5600 2.2700 ;
	    RECT 1.4200 1.8150 3.5600 1.9550 ;
	    RECT 1.4150 1.7850 3.5600 1.8150 ;
	    RECT 1.4150 1.7800 1.6650 1.7850 ;
	    RECT 1.4150 1.7750 1.6550 1.7800 ;
	    RECT 1.4150 1.7650 1.6450 1.7750 ;
	    RECT 1.4150 1.7500 1.6300 1.7650 ;
	    RECT 1.4150 1.7400 1.6250 1.7500 ;
	    RECT 1.4150 1.7250 1.6200 1.7400 ;
	    RECT 1.4150 1.7150 1.6100 1.7250 ;
	    RECT 1.4150 1.7000 1.6000 1.7150 ;
	    RECT 1.4150 1.6550 1.5850 1.7000 ;
	    RECT 1.2900 1.2450 1.5850 1.6550 ;
	    RECT 0.0850 0.9200 0.7650 1.1300 ;
	    RECT 1.4150 1.1300 1.5850 1.2450 ;
	    RECT 1.4150 0.9200 3.0550 1.1300 ;
	    RECT 0.0850 0.4050 0.3500 0.9200 ;
	    RECT 1.9850 0.3800 2.1550 0.9200 ;
	    RECT 2.8850 0.3800 3.0550 0.9200 ;
   END
END efs8hd_or4b_2
MACRO efs8hd_or4bb_2
   CLASS CORE ;
   FOREIGN efs8hd_or4bb_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 4.6000 BY 3.4000 ;
   SITE unitehd ;
   PIN CN
      PORT
         LAYER li1 ;
	    RECT 0.4300 1.1050 0.7800 2.1200 ;
      END
   END CN
   PIN DN
      PORT
         LAYER li1 ;
	    RECT 0.9500 1.1050 1.2400 1.6550 ;
      END
   END DN
   PIN A
      PORT
         LAYER li1 ;
	    RECT 2.6400 1.1050 3.2950 1.6550 ;
      END
   END A
   PIN X
      PORT
         LAYER li1 ;
	    RECT 3.8050 1.8700 4.0800 3.0800 ;
	    RECT 3.9100 0.9500 4.0800 1.8700 ;
	    RECT 3.8050 0.5200 4.0800 0.9500 ;
      END
   END X
   PIN B
      PORT
         LAYER li1 ;
	    RECT 2.4450 2.4650 3.1450 3.0700 ;
      END
   END B
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.6600 0.1050 0.8300 0.9350 ;
	    RECT 1.4950 0.1050 1.8500 0.5950 ;
	    RECT 2.3950 0.1050 2.7250 0.5950 ;
	    RECT 3.2350 0.1050 3.6150 0.5950 ;
	    RECT 4.2500 0.1050 4.4200 1.2800 ;
	    RECT 0.6600 0.0850 4.4200 0.1050 ;
	    RECT 0.0000 -0.0850 4.6000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 4.6000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 4.6000 3.4850 ;
	    RECT 0.5150 3.2950 4.4200 3.3150 ;
	    RECT 0.5150 2.7550 0.8450 3.2950 ;
	    RECT 3.3150 2.2950 3.5950 3.2950 ;
	    RECT 4.2500 1.8000 4.4200 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 4.6000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.5450 0.3450 3.0700 ;
	    RECT 1.5350 2.7550 2.2750 2.9700 ;
	    RECT 0.0850 2.3300 1.9350 2.5450 ;
	    RECT 0.0850 0.9350 0.2600 2.3300 ;
	    RECT 0.9950 1.9050 1.5950 2.1200 ;
	    RECT 1.4100 1.5550 1.5950 1.9050 ;
	    RECT 1.7650 1.9550 1.9350 2.3300 ;
	    RECT 2.1050 2.2950 2.2750 2.7550 ;
	    RECT 2.1050 2.1250 3.1450 2.2950 ;
	    RECT 2.9750 2.0800 3.1450 2.1250 ;
	    RECT 1.7650 1.7700 2.4200 1.9550 ;
	    RECT 2.9750 1.8700 3.6350 2.0800 ;
	    RECT 1.4100 1.3450 1.8550 1.5550 ;
	    RECT 1.4100 0.9350 1.6000 1.3450 ;
	    RECT 2.2500 1.2450 2.4200 1.7700 ;
	    RECT 3.4650 1.6550 3.6350 1.8700 ;
	    RECT 3.4650 1.2450 3.7400 1.6550 ;
	    RECT 3.4650 0.9350 3.6350 1.2450 ;
	    RECT 0.0850 0.5650 0.4650 0.9350 ;
	    RECT 1.0800 0.7650 1.6000 0.9350 ;
	    RECT 2.0250 0.7650 3.6350 0.9350 ;
	    RECT 1.0800 0.5650 1.2500 0.7650 ;
	    RECT 2.0250 0.3800 2.1950 0.7650 ;
	    RECT 2.8950 0.3800 3.0650 0.7650 ;
   END
END efs8hd_or4bb_2
MACRO efs8hd_sdfbbn_2
   CLASS CORE ;
   FOREIGN efs8hd_sdfbbn_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 15.1800 BY 3.4000 ;
   SITE unitehd ;
   PIN SCD
      PORT
         LAYER li1 ;
	    RECT 1.4150 1.2800 1.6950 2.1050 ;
      END
   END SCD
   PIN SCE
      PORT
         LAYER li1 ;
	    RECT 1.9350 1.3700 2.1550 2.1200 ;
	    RECT 1.9350 0.9550 2.3350 1.3700 ;
	    RECT 1.9350 0.4300 2.1450 0.9550 ;
      END
   END SCE
   PIN RESETB
      PORT
         LAYER li1 ;
	    RECT 11.5900 1.3700 12.0700 1.6550 ;
      END
   END RESETB
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.4300 0.1050 1.7050 0.7950 ;
	    RECT 3.3700 0.1050 3.7000 0.5550 ;
	    RECT 5.8850 0.1050 6.0550 0.6550 ;
	    RECT 7.6450 0.1050 7.9750 0.5800 ;
	    RECT 9.5600 0.1050 9.8200 0.6550 ;
	    RECT 12.0800 0.1050 12.4100 1.0050 ;
	    RECT 13.0000 0.1050 13.2350 1.1050 ;
	    RECT 13.9500 0.1050 14.2450 0.6800 ;
	    RECT 14.8350 0.1050 15.0750 1.1050 ;
	    RECT 0.0000 -0.1050 15.1800 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 15.1800 0.3000 ;
      END
   END vgnd
   PIN CLKN
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.2200 0.4350 2.0300 ;
      END
   END CLKN
   PIN SETB
      PORT
         LAYER li1 ;
	    RECT 5.8850 1.2050 6.2150 1.3300 ;
	    RECT 5.8850 0.9200 6.2950 1.2050 ;
	    RECT 9.7550 0.9200 10.1300 1.3300 ;
         LAYER met1 ;
	    RECT 6.0650 1.1500 6.3550 1.2050 ;
	    RECT 9.7450 1.1500 10.0350 1.2050 ;
	    RECT 6.0650 0.9750 10.0350 1.1500 ;
	    RECT 6.0650 0.9200 6.3550 0.9750 ;
	    RECT 9.7450 0.9200 10.0350 0.9750 ;
      END
   END SETB
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 14.4150 1.8050 14.6650 3.0800 ;
	    RECT 14.4600 1.0300 14.6650 1.8050 ;
	    RECT 14.4150 0.3200 14.6650 1.0300 ;
      END
   END Q
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 15.1800 3.5050 ;
	    RECT 0.5150 2.6700 0.8450 3.2950 ;
	    RECT 1.4300 2.3550 1.7850 3.2950 ;
	    RECT 3.2950 2.7700 3.6400 3.2950 ;
	    RECT 5.7050 2.7550 6.0850 3.2950 ;
	    RECT 7.1750 2.3950 7.5050 3.2950 ;
	    RECT 9.6200 2.8200 10.0000 3.2950 ;
	    RECT 10.9400 2.8200 12.4100 3.2950 ;
	    RECT 13.0000 1.8700 13.2350 3.2950 ;
	    RECT 13.9500 2.2050 14.2450 3.2950 ;
	    RECT 14.8350 1.8700 15.0750 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 15.1800 3.7000 ;
      END
   END vpwr
   PIN D
      PORT
         LAYER li1 ;
	    RECT 3.8250 1.6550 4.0250 2.9700 ;
      END
   END D
   PIN QN
      PORT
         LAYER li1 ;
	    RECT 12.5800 2.0400 12.8300 3.0800 ;
	    RECT 12.6600 0.8950 12.8300 2.0400 ;
	    RECT 12.5800 0.3200 12.8300 0.8950 ;
      END
   END QN
   OBS
         LAYER li1 ;
	    RECT 0.1700 2.4550 0.3450 3.0800 ;
	    RECT 0.1700 2.2450 0.8350 2.4550 ;
	    RECT 0.6050 1.0050 0.8350 2.2450 ;
	    RECT 0.1700 0.7950 0.8350 1.0050 ;
	    RECT 0.1700 0.4300 0.3450 0.7950 ;
	    RECT 1.0150 0.4300 1.2350 3.0800 ;
	    RECT 2.2150 2.3450 2.5750 2.9800 ;
	    RECT 2.8950 2.3800 3.0650 3.0800 ;
	    RECT 2.4050 1.7550 2.5750 2.3450 ;
	    RECT 2.7450 2.1800 3.0650 2.3800 ;
	    RECT 2.7450 1.9700 3.6450 2.1800 ;
	    RECT 2.4050 1.5650 3.0750 1.7550 ;
	    RECT 2.4350 1.5450 3.0750 1.5650 ;
	    RECT 2.5600 1.3450 3.0750 1.5450 ;
	    RECT 3.4750 1.3700 3.6450 1.9700 ;
	    RECT 2.5600 0.7450 2.7300 1.3450 ;
	    RECT 3.4750 0.9950 3.7700 1.3700 ;
	    RECT 2.3150 0.3300 2.7300 0.7450 ;
	    RECT 2.9550 0.9550 3.7700 0.9950 ;
	    RECT 2.9550 0.7800 3.6450 0.9550 ;
	    RECT 2.9550 0.3800 3.1250 0.7800 ;
	    RECT 4.2300 0.3800 4.4550 3.0800 ;
	    RECT 4.6350 2.8150 5.4650 3.0250 ;
	    RECT 4.6250 1.9700 5.1250 2.4450 ;
	    RECT 4.6250 0.8800 4.8450 1.9700 ;
	    RECT 5.2950 1.7550 5.4650 2.8150 ;
	    RECT 6.3850 2.5450 6.5550 2.9700 ;
	    RECT 8.5500 2.8150 9.3800 3.0250 ;
	    RECT 5.6350 2.2300 6.9850 2.5450 ;
	    RECT 5.6350 1.9700 5.8850 2.2300 ;
	    RECT 6.3950 1.7550 6.6450 1.8550 ;
	    RECT 5.2950 1.5450 6.6450 1.7550 ;
	    RECT 5.2950 1.4950 5.7150 1.5450 ;
	    RECT 5.0250 0.8050 5.3750 1.2700 ;
	    RECT 5.5450 0.5800 5.7150 1.4950 ;
	    RECT 6.4250 1.4450 6.6450 1.5450 ;
	    RECT 6.8150 1.3300 6.9850 2.2300 ;
	    RECT 7.1550 1.7700 8.1600 2.0700 ;
	    RECT 8.3600 1.9700 8.5950 2.4800 ;
	    RECT 7.1550 1.5450 7.4850 1.7700 ;
	    RECT 8.8350 1.6300 9.0400 2.3800 ;
	    RECT 7.7950 1.3300 8.1250 1.5450 ;
	    RECT 6.8150 1.1200 8.1250 1.3300 ;
	    RECT 8.4200 1.4050 9.0400 1.6300 ;
	    RECT 9.2100 1.7550 9.3800 2.8150 ;
	    RECT 10.2400 2.6050 10.4100 2.9700 ;
	    RECT 9.5500 2.3950 12.4100 2.6050 ;
	    RECT 9.5500 1.9700 9.8000 2.3950 ;
	    RECT 9.2100 1.5450 10.5600 1.7550 ;
	    RECT 6.8150 0.9550 7.0350 1.1200 ;
	    RECT 6.7050 0.7450 7.0350 0.9550 ;
	    RECT 4.7000 0.3300 5.7150 0.5800 ;
	    RECT 6.2250 0.5300 6.5550 0.6300 ;
	    RECT 7.2050 0.5300 7.3750 0.8950 ;
	    RECT 8.4200 0.8800 8.7050 1.4050 ;
	    RECT 9.2100 0.5800 9.3800 1.5450 ;
	    RECT 10.3400 1.3450 10.5600 1.5450 ;
	    RECT 10.7300 0.9750 10.9100 2.3950 ;
	    RECT 10.5800 0.7450 10.9100 0.9750 ;
	    RECT 11.0800 1.9700 11.9250 2.1800 ;
	    RECT 11.0800 1.1550 11.3550 1.9700 ;
	    RECT 12.2400 1.6550 12.4100 2.3950 ;
	    RECT 13.4550 1.6550 13.7700 3.0200 ;
	    RECT 12.2400 1.2450 12.4800 1.6550 ;
	    RECT 13.4550 1.2450 14.2900 1.6550 ;
	    RECT 11.0800 0.9450 11.8450 1.1550 ;
	    RECT 6.2250 0.3200 7.3750 0.5300 ;
	    RECT 8.6150 0.3300 9.3800 0.5800 ;
	    RECT 10.0800 0.5300 10.4100 0.6800 ;
	    RECT 11.0800 0.5300 11.2500 0.7300 ;
	    RECT 10.0800 0.3200 11.2500 0.5300 ;
	    RECT 11.6200 0.3300 11.8450 0.9450 ;
	    RECT 13.4550 0.3200 13.7700 1.2450 ;
         LAYER met1 ;
	    RECT 1.0050 2.4250 1.2950 2.4800 ;
	    RECT 4.6850 2.4250 4.9750 2.4800 ;
	    RECT 8.3650 2.4250 8.6550 2.4800 ;
	    RECT 1.0050 2.2500 8.6550 2.4250 ;
	    RECT 1.0050 2.1950 1.2950 2.2500 ;
	    RECT 4.6850 2.1950 4.9750 2.2500 ;
	    RECT 8.3650 2.1950 8.6550 2.2500 ;
	    RECT 7.9050 2.0000 8.1950 2.0550 ;
	    RECT 11.1250 2.0000 11.4150 2.0550 ;
	    RECT 7.9050 1.8250 11.4150 2.0000 ;
	    RECT 7.9050 1.7700 8.1950 1.8250 ;
	    RECT 11.1250 1.7700 11.4150 1.8250 ;
	    RECT 2.8450 1.5750 3.1350 1.6300 ;
	    RECT 4.2250 1.5750 4.5150 1.6300 ;
	    RECT 8.3650 1.5750 8.6550 1.6300 ;
	    RECT 2.8450 1.4000 4.5150 1.5750 ;
	    RECT 2.8450 1.3450 3.1350 1.4000 ;
	    RECT 4.2250 1.3450 4.5150 1.4000 ;
	    RECT 5.2200 1.4000 8.6550 1.5750 ;
	    RECT 5.2200 1.2050 5.4350 1.4000 ;
	    RECT 8.3650 1.3450 8.6550 1.4000 ;
	    RECT 0.5450 1.1500 0.8350 1.2050 ;
	    RECT 5.1450 1.1500 5.4350 1.2050 ;
	    RECT 0.5450 0.9750 5.4350 1.1500 ;
	    RECT 0.5450 0.9200 0.8350 0.9750 ;
	    RECT 5.1450 0.9200 5.4350 0.9750 ;
   END
END efs8hd_sdfbbn_2
MACRO efs8hd_sdfrbp_2
   CLASS CORE ;
   FOREIGN efs8hd_sdfrbp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 13.3400 BY 3.4000 ;
   SITE unitehd ;
   PIN RESETB
      PORT
         LAYER li1 ;
	    RECT 9.5250 1.3300 10.1150 1.6150 ;
	    RECT 6.5050 0.9550 7.0350 1.3050 ;
	    RECT 9.8050 0.7650 10.1150 1.3300 ;
         LAYER met1 ;
	    RECT 9.6300 1.2050 9.9200 1.6300 ;
	    RECT 6.4450 1.1500 7.0950 1.2050 ;
	    RECT 9.6300 1.1500 10.1750 1.2050 ;
	    RECT 6.4450 0.9750 10.1750 1.1500 ;
	    RECT 6.4450 0.9200 7.0950 0.9750 ;
	    RECT 9.8850 0.9200 10.1750 0.9750 ;
      END
   END RESETB
   PIN QN
      PORT
         LAYER li1 ;
	    RECT 12.5250 2.6000 12.8250 3.0800 ;
	    RECT 12.4350 1.9200 12.8250 2.6000 ;
	    RECT 12.6550 1.0300 12.8250 1.9200 ;
	    RECT 12.4450 0.3900 12.8250 1.0300 ;
      END
   END QN
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 11.5750 0.3300 11.9250 2.1200 ;
      END
   END Q
   PIN CLK
      PORT
         LAYER li1 ;
	    RECT 0.1400 1.1050 0.4900 2.0300 ;
      END
   END CLK
   PIN SCE
      PORT
         LAYER li1 ;
	    RECT 1.4650 2.4800 1.7300 3.0800 ;
	    RECT 1.4850 1.3400 1.7300 2.4800 ;
      END
   END SCE
   PIN D
      PORT
         LAYER li1 ;
	    RECT 2.8650 2.2300 3.1200 3.0800 ;
	    RECT 2.7350 1.6950 3.1200 2.2300 ;
      END
   END D
   PIN SCD
      PORT
         LAYER li1 ;
	    RECT 4.0200 0.8900 4.4550 2.1250 ;
	    RECT 4.0200 0.3550 4.2750 0.8900 ;
      END
   END SCD
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.8750 0.1050 2.2050 0.7000 ;
	    RECT 2.3950 0.1050 2.7250 1.0300 ;
	    RECT 4.4450 0.1050 4.7750 0.6750 ;
	    RECT 6.9150 0.1050 7.2450 0.6800 ;
	    RECT 9.0850 0.1050 9.2550 0.6550 ;
	    RECT 11.0900 0.1050 11.3650 0.6800 ;
	    RECT 12.1050 0.1050 12.2750 1.0300 ;
	    RECT 12.9950 0.1050 13.1650 1.1650 ;
	    RECT 0.5150 0.0850 13.1650 0.1050 ;
	    RECT 0.0000 -0.0850 13.3400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 13.3400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 13.3400 3.4850 ;
	    RECT 0.5300 3.2950 13.2450 3.3150 ;
	    RECT 0.5300 2.6700 0.8600 3.2950 ;
	    RECT 2.3200 2.5500 2.4900 3.2950 ;
	    RECT 4.3000 2.8450 4.6300 3.2950 ;
	    RECT 6.4100 2.9450 6.7400 3.2950 ;
	    RECT 7.3750 2.7200 7.7450 3.2950 ;
	    RECT 9.3600 2.7450 9.6100 3.2950 ;
	    RECT 10.1200 2.8200 10.4500 3.2950 ;
	    RECT 11.0900 2.7550 11.4200 3.2950 ;
	    RECT 12.0250 2.8200 12.3550 3.2950 ;
	    RECT 12.9950 1.8700 13.2450 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 13.3400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0900 2.4550 0.3450 3.0800 ;
	    RECT 0.0900 2.2450 0.8650 2.4550 ;
	    RECT 0.6600 1.6550 0.8650 2.2450 ;
	    RECT 1.0350 2.3750 1.2050 3.0800 ;
	    RECT 1.9000 2.5700 2.1500 3.0000 ;
	    RECT 3.4600 2.6300 3.6300 3.0800 ;
	    RECT 4.9050 2.7300 5.2750 3.0450 ;
	    RECT 4.9050 2.6300 5.0750 2.7300 ;
	    RECT 5.4700 2.6700 5.8350 3.0800 ;
	    RECT 1.0350 2.1650 1.3150 2.3750 ;
	    RECT 0.6600 1.2450 0.9750 1.6550 ;
	    RECT 0.6600 0.9350 0.8350 1.2450 ;
	    RECT 0.0950 0.7650 0.8350 0.9350 ;
	    RECT 1.1450 0.8450 1.3150 2.1650 ;
	    RECT 1.9800 1.8200 2.1500 2.5700 ;
	    RECT 3.2900 2.4200 5.0750 2.6300 ;
	    RECT 1.9800 1.5750 2.4700 1.8200 ;
	    RECT 2.0550 1.4800 2.4700 1.5750 ;
	    RECT 3.2900 1.4800 3.4600 2.4200 ;
	    RECT 2.0550 1.2450 3.0850 1.4800 ;
	    RECT 2.0550 1.1250 2.2250 1.2450 ;
	    RECT 0.0950 0.4300 0.3450 0.7650 ;
	    RECT 1.0150 0.4300 1.3150 0.8450 ;
	    RECT 1.5350 0.9150 2.2250 1.1250 ;
	    RECT 1.5350 0.4950 1.7050 0.9150 ;
	    RECT 2.9150 0.5300 3.0850 1.2450 ;
	    RECT 3.2550 1.2700 3.4600 1.4800 ;
	    RECT 3.2550 0.8450 3.4250 1.2700 ;
	    RECT 3.6800 0.5300 3.8500 2.1050 ;
	    RECT 4.6250 1.1200 4.7950 2.4200 ;
	    RECT 5.2450 1.9700 5.4950 2.4450 ;
	    RECT 4.9650 1.3300 5.1350 1.7450 ;
	    RECT 5.3250 1.2950 5.4950 1.9700 ;
	    RECT 5.6650 1.7300 5.8350 2.6700 ;
	    RECT 6.0050 2.6300 6.1750 2.9700 ;
	    RECT 6.9950 2.6300 7.1650 2.9700 ;
	    RECT 6.0050 2.4200 7.1650 2.6300 ;
	    RECT 7.9700 2.5050 8.1400 3.0800 ;
	    RECT 8.3200 2.6550 9.1900 3.0800 ;
	    RECT 9.0150 2.6450 9.1900 2.6550 ;
	    RECT 9.0150 2.5450 9.2100 2.6450 ;
	    RECT 7.4550 2.2950 8.1400 2.5050 ;
	    RECT 8.3100 2.4200 8.8400 2.4450 ;
	    RECT 7.4550 2.2050 7.7150 2.2950 ;
	    RECT 6.2850 1.9950 7.7150 2.2050 ;
	    RECT 8.3100 2.0800 8.8700 2.4200 ;
	    RECT 5.6650 1.5200 7.3750 1.7300 ;
	    RECT 4.6250 0.8950 5.1450 1.1200 ;
	    RECT 2.9150 0.3200 3.8500 0.5300 ;
	    RECT 4.9750 0.6300 5.1450 0.8950 ;
	    RECT 5.3250 0.8800 5.9750 1.2950 ;
	    RECT 4.9750 0.4200 5.3150 0.6300 ;
	    RECT 6.1650 0.5950 6.3350 1.5200 ;
	    RECT 7.2050 1.2550 7.3750 1.5200 ;
	    RECT 7.5450 1.0450 7.7150 1.9950 ;
	    RECT 5.4850 0.3800 6.3350 0.5950 ;
	    RECT 7.4550 0.5550 7.7150 1.0450 ;
	    RECT 7.8850 2.0700 8.8700 2.0800 ;
	    RECT 9.0400 2.1800 9.2100 2.5450 ;
	    RECT 9.7800 2.6050 9.9500 2.9700 ;
	    RECT 9.7800 2.3950 10.5450 2.6050 ;
	    RECT 7.8850 1.8700 8.5200 2.0700 ;
	    RECT 9.0400 1.9700 10.2050 2.1800 ;
	    RECT 7.8850 0.8800 8.0950 1.8700 ;
	    RECT 9.0400 1.8550 9.2100 1.9700 ;
	    RECT 8.4050 1.1500 8.5750 1.6550 ;
	    RECT 8.7450 1.6450 9.2100 1.8550 ;
	    RECT 10.3750 1.6550 10.5450 2.3950 ;
	    RECT 10.7150 2.5450 10.8900 3.0800 ;
	    RECT 11.5500 2.5450 12.2650 2.6050 ;
	    RECT 10.7150 2.3300 12.2650 2.5450 ;
	    RECT 10.7150 2.2450 11.4050 2.3300 ;
	    RECT 8.7450 0.6700 8.9150 1.6450 ;
	    RECT 10.3750 1.6200 11.0600 1.6550 ;
	    RECT 9.1250 1.0800 9.2950 1.4300 ;
	    RECT 10.3450 1.3200 11.0600 1.6200 ;
	    RECT 9.1250 0.8700 9.6350 1.0800 ;
	    RECT 7.4550 0.3450 7.7850 0.5550 ;
	    RECT 8.0050 0.3200 8.9150 0.6700 ;
	    RECT 9.4650 0.5800 9.6350 0.8700 ;
	    RECT 10.3450 0.5800 10.5150 1.3200 ;
	    RECT 11.2300 1.1050 11.4050 2.2450 ;
	    RECT 12.0950 1.6550 12.2650 2.3300 ;
	    RECT 12.0950 1.2450 12.4850 1.6550 ;
	    RECT 9.4650 0.3700 10.5150 0.5800 ;
	    RECT 10.7150 0.8950 11.4050 1.1050 ;
	    RECT 10.7150 0.4300 10.8850 0.8950 ;
         LAYER met1 ;
	    RECT 0.9700 2.4250 1.2700 2.4800 ;
	    RECT 5.2650 2.4250 5.5550 2.4800 ;
	    RECT 8.3850 2.4250 8.6750 2.4800 ;
	    RECT 0.9700 2.2500 8.6750 2.4250 ;
	    RECT 0.9700 2.1950 1.2700 2.2500 ;
	    RECT 5.2650 2.1950 5.5550 2.2500 ;
	    RECT 8.3850 2.1950 8.6750 2.2500 ;
	    RECT 0.7450 1.5750 1.0350 1.6300 ;
	    RECT 4.8450 1.5800 5.1350 1.6300 ;
	    RECT 8.3450 1.5800 8.6350 1.6300 ;
	    RECT 4.8450 1.5750 8.6350 1.5800 ;
	    RECT 0.7450 1.4000 8.6350 1.5750 ;
	    RECT 0.7450 1.3450 1.0350 1.4000 ;
	    RECT 4.8450 1.3500 8.6350 1.4000 ;
	    RECT 4.8450 1.3450 5.1350 1.3500 ;
	    RECT 8.3450 1.3450 8.6350 1.3500 ;
   END
END efs8hd_sdfrbp_2
MACRO efs8hd_sdfrtp_2
   CLASS CORE ;
   FOREIGN efs8hd_sdfrtp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 11.9600 BY 3.4000 ;
   SITE unitehd ;
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 11.1400 1.8250 11.4000 2.9050 ;
	    RECT 11.1500 1.8050 11.4000 1.8250 ;
	    RECT 11.1900 0.9950 11.4000 1.8050 ;
	    RECT 11.1400 0.3300 11.4000 0.9950 ;
      END
   END Q
   PIN RESETB
      PORT
         LAYER li1 ;
	    RECT 9.5250 1.3300 10.1150 1.6150 ;
	    RECT 6.5050 0.9550 7.0350 1.3050 ;
	    RECT 9.8050 0.7650 10.1150 1.3300 ;
         LAYER met1 ;
	    RECT 9.6300 1.2050 9.9200 1.6300 ;
	    RECT 6.4450 1.1500 7.0950 1.2050 ;
	    RECT 9.6300 1.1500 10.1750 1.2050 ;
	    RECT 6.4450 0.9750 10.1750 1.1500 ;
	    RECT 6.4450 0.9200 7.0950 0.9750 ;
	    RECT 9.8850 0.9200 10.1750 0.9750 ;
      END
   END RESETB
   PIN CLK
      PORT
         LAYER li1 ;
	    RECT 0.1400 1.1050 0.4900 2.0300 ;
      END
   END CLK
   PIN SCE
      PORT
         LAYER li1 ;
	    RECT 1.4650 2.4800 1.7300 3.0800 ;
	    RECT 1.4850 1.3400 1.7300 2.4800 ;
      END
   END SCE
   PIN D
      PORT
         LAYER li1 ;
	    RECT 2.8650 2.2300 3.1200 3.0800 ;
	    RECT 2.7350 1.6950 3.1200 2.2300 ;
      END
   END D
   PIN SCD
      PORT
         LAYER li1 ;
	    RECT 4.0200 0.8900 4.4550 2.1250 ;
	    RECT 4.0200 0.3550 4.2750 0.8900 ;
      END
   END SCD
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.8750 0.1050 2.2050 0.7000 ;
	    RECT 2.3950 0.1050 2.7250 1.0300 ;
	    RECT 4.4450 0.1050 4.7750 0.6750 ;
	    RECT 6.9150 0.1050 7.2450 0.6800 ;
	    RECT 9.0850 0.1050 9.2550 0.6550 ;
	    RECT 10.7200 0.1050 10.8900 0.6800 ;
	    RECT 11.5700 0.1050 11.7400 0.6800 ;
	    RECT 0.5150 0.0850 11.7400 0.1050 ;
	    RECT 0.0000 -0.0850 11.9600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 11.9600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 11.9600 3.4850 ;
	    RECT 0.5300 3.2950 11.8200 3.3150 ;
	    RECT 0.5300 2.6700 0.8600 3.2950 ;
	    RECT 2.3200 2.5500 2.4900 3.2950 ;
	    RECT 4.3000 2.8450 4.6300 3.2950 ;
	    RECT 6.4100 2.9450 6.7400 3.2950 ;
	    RECT 7.3750 2.7200 7.7450 3.2950 ;
	    RECT 9.3600 2.7450 9.6100 3.2950 ;
	    RECT 10.1200 2.8200 10.4500 3.2950 ;
	    RECT 10.7200 1.8700 10.9700 3.2950 ;
	    RECT 11.5700 1.8700 11.8200 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 11.9600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0900 2.4550 0.3450 3.0800 ;
	    RECT 0.0900 2.2450 0.8650 2.4550 ;
	    RECT 0.6600 1.6550 0.8650 2.2450 ;
	    RECT 1.0350 2.3750 1.2050 3.0800 ;
	    RECT 1.9000 2.5700 2.1500 3.0000 ;
	    RECT 3.4600 2.6300 3.6300 3.0800 ;
	    RECT 4.9050 2.7300 5.2750 3.0450 ;
	    RECT 4.9050 2.6300 5.0750 2.7300 ;
	    RECT 5.4700 2.6700 5.8350 3.0800 ;
	    RECT 1.0350 2.1650 1.3150 2.3750 ;
	    RECT 0.6600 1.2450 0.9750 1.6550 ;
	    RECT 0.6600 0.9350 0.8350 1.2450 ;
	    RECT 0.0950 0.7650 0.8350 0.9350 ;
	    RECT 1.1450 0.8450 1.3150 2.1650 ;
	    RECT 1.9800 1.8200 2.1500 2.5700 ;
	    RECT 3.2900 2.4200 5.0750 2.6300 ;
	    RECT 1.9800 1.5750 2.4700 1.8200 ;
	    RECT 2.0550 1.4800 2.4700 1.5750 ;
	    RECT 3.2900 1.4800 3.4600 2.4200 ;
	    RECT 2.0550 1.2450 3.0850 1.4800 ;
	    RECT 2.0550 1.1250 2.2250 1.2450 ;
	    RECT 0.0950 0.4300 0.3450 0.7650 ;
	    RECT 1.0150 0.4300 1.3150 0.8450 ;
	    RECT 1.5350 0.9150 2.2250 1.1250 ;
	    RECT 1.5350 0.4950 1.7050 0.9150 ;
	    RECT 2.9150 0.5300 3.0850 1.2450 ;
	    RECT 3.2550 1.2700 3.4600 1.4800 ;
	    RECT 3.2550 0.8450 3.4250 1.2700 ;
	    RECT 3.6800 0.5300 3.8500 2.1050 ;
	    RECT 4.6250 1.1200 4.7950 2.4200 ;
	    RECT 5.2450 1.9700 5.4950 2.4450 ;
	    RECT 4.9650 1.3300 5.1350 1.7450 ;
	    RECT 5.3250 1.2950 5.4950 1.9700 ;
	    RECT 5.6650 1.7300 5.8350 2.6700 ;
	    RECT 6.0050 2.6300 6.1750 2.9700 ;
	    RECT 6.9950 2.6300 7.1650 2.9700 ;
	    RECT 6.0050 2.4200 7.1650 2.6300 ;
	    RECT 7.9700 2.5050 8.1400 3.0800 ;
	    RECT 8.3200 2.6550 9.1900 3.0800 ;
	    RECT 9.0150 2.6450 9.1900 2.6550 ;
	    RECT 9.0150 2.5450 9.2100 2.6450 ;
	    RECT 7.4550 2.2950 8.1400 2.5050 ;
	    RECT 8.3100 2.4200 8.8400 2.4450 ;
	    RECT 7.4550 2.2050 7.7150 2.2950 ;
	    RECT 6.2850 1.9950 7.7150 2.2050 ;
	    RECT 8.3100 2.0800 8.8700 2.4200 ;
	    RECT 5.6650 1.5200 7.3750 1.7300 ;
	    RECT 4.6250 0.8950 5.1450 1.1200 ;
	    RECT 2.9150 0.3200 3.8500 0.5300 ;
	    RECT 4.9750 0.6300 5.1450 0.8950 ;
	    RECT 5.3250 0.8800 5.9750 1.2950 ;
	    RECT 4.9750 0.4200 5.3150 0.6300 ;
	    RECT 6.1650 0.5950 6.3350 1.5200 ;
	    RECT 7.2050 1.2550 7.3750 1.5200 ;
	    RECT 7.5450 1.0450 7.7150 1.9950 ;
	    RECT 5.4850 0.3800 6.3350 0.5950 ;
	    RECT 7.4550 0.5550 7.7150 1.0450 ;
	    RECT 7.8850 2.0700 8.8700 2.0800 ;
	    RECT 9.0400 2.1800 9.2100 2.5450 ;
	    RECT 9.7800 2.6050 9.9500 2.9700 ;
	    RECT 9.7800 2.3950 10.5450 2.6050 ;
	    RECT 7.8850 1.8700 8.5200 2.0700 ;
	    RECT 9.0400 1.9700 10.2050 2.1800 ;
	    RECT 7.8850 0.8800 8.0950 1.8700 ;
	    RECT 9.0400 1.8550 9.2100 1.9700 ;
	    RECT 8.4050 1.1500 8.5750 1.6550 ;
	    RECT 8.7450 1.6450 9.2100 1.8550 ;
	    RECT 10.3750 1.6550 10.5450 2.3950 ;
	    RECT 8.7450 0.6700 8.9150 1.6450 ;
	    RECT 10.3750 1.6200 11.0200 1.6550 ;
	    RECT 9.1250 1.0800 9.2950 1.4300 ;
	    RECT 10.3450 1.2450 11.0200 1.6200 ;
	    RECT 9.1250 0.8700 9.6350 1.0800 ;
	    RECT 7.4550 0.3450 7.7850 0.5550 ;
	    RECT 8.0050 0.3200 8.9150 0.6700 ;
	    RECT 9.4650 0.5800 9.6350 0.8700 ;
	    RECT 10.3450 0.5800 10.5150 1.2450 ;
	    RECT 9.4650 0.3700 10.5150 0.5800 ;
         LAYER met1 ;
	    RECT 0.9700 2.4250 1.2700 2.4800 ;
	    RECT 5.2650 2.4250 5.5550 2.4800 ;
	    RECT 8.3850 2.4250 8.6750 2.4800 ;
	    RECT 0.9700 2.2500 8.6750 2.4250 ;
	    RECT 0.9700 2.1950 1.2700 2.2500 ;
	    RECT 5.2650 2.1950 5.5550 2.2500 ;
	    RECT 8.3850 2.1950 8.6750 2.2500 ;
	    RECT 0.7450 1.5750 1.0350 1.6300 ;
	    RECT 4.8450 1.6050 5.1350 1.6300 ;
	    RECT 8.3450 1.6050 8.6350 1.6300 ;
	    RECT 4.8450 1.5750 8.6350 1.6050 ;
	    RECT 0.7450 1.4000 8.6350 1.5750 ;
	    RECT 0.7450 1.3450 1.0350 1.4000 ;
	    RECT 4.8450 1.3750 8.6350 1.4000 ;
	    RECT 4.8450 1.3450 5.1350 1.3750 ;
	    RECT 8.3450 1.3450 8.6350 1.3750 ;
   END
END efs8hd_sdfrtp_2
MACRO efs8hd_sdfsbp_2
   CLASS CORE ;
   FOREIGN efs8hd_sdfsbp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 14.2600 BY 3.4000 ;
   SITE unitehd ;
   PIN QN
      PORT
         LAYER li1 ;
	    RECT 11.4600 0.3200 11.8550 3.0800 ;
      END
   END QN
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 13.4100 1.8700 13.7400 3.0650 ;
	    RECT 13.5150 1.0300 13.7400 1.8700 ;
	    RECT 13.4100 0.3450 13.7400 1.0300 ;
      END
   END Q
   PIN SCD
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.9550 0.3400 2.0950 ;
      END
   END SCD
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.0500 0.9550 1.3350 2.0950 ;
      END
   END D
   PIN CLK
      PORT
         LAYER li1 ;
	    RECT 2.9050 2.0200 3.1000 2.4650 ;
	    RECT 2.9050 1.3200 3.5650 2.0200 ;
	    RECT 2.9050 0.9050 3.1000 1.3200 ;
      END
   END CLK
   PIN SCE
      PORT
         LAYER li1 ;
	    RECT 0.5400 0.9550 0.8200 2.0950 ;
	    RECT 2.4050 1.3450 2.7350 1.9900 ;
         LAYER met1 ;
	    RECT 0.5450 1.5750 0.8350 1.6300 ;
	    RECT 2.3850 1.5750 2.6750 1.6300 ;
	    RECT 0.5450 1.4000 2.6750 1.5750 ;
	    RECT 0.5450 1.3450 0.8350 1.4000 ;
	    RECT 2.3850 1.3450 2.6750 1.4000 ;
      END
   END SCE
   PIN SETB
      PORT
         LAYER li1 ;
	    RECT 6.5850 1.7850 7.0650 2.2950 ;
	    RECT 8.8800 1.9050 9.9350 2.1550 ;
	    RECT 8.8800 1.7950 9.1150 1.9050 ;
         LAYER met1 ;
	    RECT 6.5800 2.0000 6.8700 2.0550 ;
	    RECT 8.8800 2.0000 9.1700 2.0550 ;
	    RECT 6.5800 1.8250 9.1700 2.0000 ;
	    RECT 6.5800 1.7700 6.8700 1.8250 ;
	    RECT 8.8800 1.7700 9.1700 1.8250 ;
      END
   END SETB
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.1050 0.7000 0.7450 ;
	    RECT 1.8400 0.1050 2.0900 0.6800 ;
	    RECT 2.7000 0.1050 3.1000 0.6950 ;
	    RECT 3.6400 0.1050 3.9400 0.6800 ;
	    RECT 5.6650 0.1050 6.1650 0.5800 ;
	    RECT 6.7200 0.1050 7.7050 1.0050 ;
	    RECT 10.0350 0.1050 10.2850 0.6800 ;
	    RECT 11.1200 0.1050 11.2900 1.1050 ;
	    RECT 12.0250 0.1050 12.3150 1.1050 ;
	    RECT 12.8850 0.1050 13.2400 1.0300 ;
	    RECT 13.9100 0.1050 14.1750 1.1050 ;
	    RECT 0.0850 0.0850 14.1750 0.1050 ;
	    RECT 0.0000 -0.0850 14.2600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 14.2600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 14.2600 3.4850 ;
	    RECT 0.5150 3.2950 14.1750 3.3150 ;
	    RECT 0.5150 2.8450 0.8450 3.2950 ;
	    RECT 2.7050 2.6750 3.1000 3.2950 ;
	    RECT 3.6450 2.8450 3.9750 3.2950 ;
	    RECT 6.0000 2.8450 6.3300 3.2950 ;
	    RECT 7.0600 2.6550 8.0150 3.2950 ;
	    RECT 9.1600 2.7950 9.4900 3.2950 ;
	    RECT 10.1000 2.7950 10.4300 3.2950 ;
	    RECT 11.0800 1.8550 11.2900 3.2950 ;
	    RECT 12.0250 1.8550 12.3150 3.2950 ;
	    RECT 12.8850 2.0450 13.2400 3.2950 ;
	    RECT 13.9100 1.8550 14.1750 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 14.2600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.5950 0.3450 3.0800 ;
	    RECT 1.0150 2.8200 2.1050 3.0800 ;
	    RECT 1.0150 2.5950 1.1850 2.8200 ;
	    RECT 2.2750 2.6050 2.5350 3.0800 ;
	    RECT 0.0850 2.3050 1.1850 2.5950 ;
	    RECT 1.3550 2.3050 1.6950 2.6050 ;
	    RECT 1.5050 0.9000 1.6950 2.3050 ;
	    RECT 1.5000 0.8800 1.6950 0.9000 ;
	    RECT 1.9800 2.2000 2.5350 2.6050 ;
	    RECT 3.2700 2.5000 3.4750 2.9050 ;
	    RECT 4.1450 2.6700 4.4400 3.0800 ;
	    RECT 3.2700 2.2900 3.9950 2.5000 ;
	    RECT 1.9800 1.1300 2.2350 2.2000 ;
	    RECT 1.9800 0.8950 2.5300 1.1300 ;
	    RECT 3.7350 1.1050 3.9950 2.2900 ;
	    RECT 1.4950 0.8050 1.6950 0.8800 ;
	    RECT 1.4950 0.7450 1.6700 0.8050 ;
	    RECT 0.8700 0.3200 1.6700 0.7450 ;
	    RECT 2.2600 0.3200 2.5300 0.8950 ;
	    RECT 3.2700 0.8950 3.9950 1.1050 ;
	    RECT 4.1650 1.7750 4.4400 2.6700 ;
	    RECT 4.6650 2.0200 4.8900 3.0800 ;
	    RECT 5.0600 2.6700 5.8050 3.0800 ;
	    RECT 4.6650 1.9900 4.9700 2.0200 ;
	    RECT 4.7150 1.8050 4.9700 1.9900 ;
	    RECT 5.2050 1.9700 5.4650 2.4450 ;
	    RECT 4.1650 1.3650 4.4900 1.7750 ;
	    RECT 3.2700 0.3200 3.4700 0.8950 ;
	    RECT 4.1650 0.7300 4.3350 1.3650 ;
	    RECT 4.7150 1.1500 4.8850 1.8050 ;
	    RECT 5.6350 1.7450 5.8050 2.6700 ;
	    RECT 6.6050 2.6350 6.8200 3.0650 ;
	    RECT 8.1850 2.6550 8.9900 3.0750 ;
	    RECT 5.9750 2.4650 6.8200 2.6350 ;
	    RECT 8.8200 2.5800 8.9900 2.6550 ;
	    RECT 9.6600 2.5800 9.9300 3.0650 ;
	    RECT 5.9750 1.9700 6.1450 2.4650 ;
	    RECT 7.3850 2.1300 8.0550 2.4450 ;
	    RECT 5.1400 1.6550 5.8050 1.7450 ;
	    RECT 5.1400 1.6100 6.4750 1.6550 ;
	    RECT 7.3550 1.6100 7.7050 1.6550 ;
	    RECT 5.1400 1.5950 7.7050 1.6100 ;
	    RECT 4.1100 0.3200 4.3350 0.7300 ;
	    RECT 4.5050 0.3200 4.8850 1.1500 ;
	    RECT 5.0550 1.4400 7.7050 1.5950 ;
	    RECT 5.0550 0.3200 5.4500 1.4400 ;
	    RECT 5.6200 1.0050 6.0150 1.2700 ;
	    RECT 6.3050 1.2200 7.7050 1.4400 ;
	    RECT 7.8850 1.1200 8.0550 2.1300 ;
	    RECT 8.4200 1.3450 8.6500 2.3800 ;
	    RECT 8.8200 2.3700 10.4300 2.5800 ;
	    RECT 10.1050 1.9050 10.4300 2.3700 ;
	    RECT 10.6000 1.6950 10.8450 3.0800 ;
	    RECT 8.8300 1.1200 9.0850 1.5800 ;
	    RECT 5.6200 0.7950 6.5500 1.0050 ;
	    RECT 7.8850 0.8700 9.0850 1.1200 ;
	    RECT 9.2850 1.4800 10.9100 1.6950 ;
	    RECT 9.2850 1.0700 9.5150 1.4800 ;
	    RECT 9.6850 1.0550 10.5600 1.2700 ;
	    RECT 6.3350 0.3200 6.5500 0.7950 ;
	    RECT 9.6850 0.6450 9.8550 1.0550 ;
	    RECT 10.7300 0.7300 10.9100 1.4800 ;
	    RECT 8.4650 0.3450 9.8550 0.6450 ;
	    RECT 10.4650 0.3200 10.9100 0.7300 ;
	    RECT 12.5300 1.6550 12.7150 3.0800 ;
	    RECT 12.5300 1.2450 13.3450 1.6550 ;
	    RECT 12.5300 0.3200 12.7150 1.2450 ;
         LAYER met1 ;
	    RECT 3.7650 2.4250 4.0550 2.4800 ;
	    RECT 5.2000 2.4250 5.4900 2.4800 ;
	    RECT 7.5000 2.4250 7.7900 2.4800 ;
	    RECT 3.7650 2.2500 7.7900 2.4250 ;
	    RECT 3.7650 2.1950 4.0550 2.2500 ;
	    RECT 5.2000 2.1950 5.4900 2.2500 ;
	    RECT 7.5000 2.1950 7.7900 2.2500 ;
	    RECT 1.4650 2.0000 1.7550 2.0550 ;
	    RECT 4.7400 2.0000 5.0300 2.0550 ;
	    RECT 1.4650 1.8250 5.0300 2.0000 ;
	    RECT 1.4650 1.7700 1.7550 1.8250 ;
	    RECT 4.7400 1.7700 5.0300 1.8250 ;
	    RECT 4.2250 1.5750 4.5150 1.6300 ;
	    RECT 8.4200 1.5750 8.7100 1.6300 ;
	    RECT 4.2250 1.4000 8.7100 1.5750 ;
	    RECT 4.2250 1.3450 4.5150 1.4000 ;
	    RECT 8.4200 1.3450 8.7100 1.4000 ;
   END
END efs8hd_sdfsbp_2
MACRO efs8hd_sdfstp_2
   CLASS CORE ;
   FOREIGN efs8hd_sdfstp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 12.8800 BY 3.4000 ;
   SITE unitehd ;
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 12.0350 1.8700 12.3650 3.0650 ;
	    RECT 12.1450 1.0300 12.3650 1.8700 ;
	    RECT 12.0350 0.3200 12.3650 1.0300 ;
      END
   END Q
   PIN SCD
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.9550 0.3400 2.0950 ;
      END
   END SCD
   PIN D
      PORT
         LAYER li1 ;
	    RECT 1.0500 0.9550 1.3350 2.0950 ;
      END
   END D
   PIN CLK
      PORT
         LAYER li1 ;
	    RECT 2.9050 2.0200 3.0850 2.4500 ;
	    RECT 2.9050 1.3200 3.5650 2.0200 ;
	    RECT 2.9050 0.9050 3.1000 1.3200 ;
      END
   END CLK
   PIN SCE
      PORT
         LAYER li1 ;
	    RECT 0.5400 0.9550 0.8200 2.0950 ;
	    RECT 2.3700 1.3450 2.7000 2.0000 ;
         LAYER met1 ;
	    RECT 0.5450 1.5750 0.8350 1.6300 ;
	    RECT 2.3850 1.5750 2.6750 1.6300 ;
	    RECT 0.5450 1.4000 2.6750 1.5750 ;
	    RECT 0.5450 1.3450 0.8350 1.4000 ;
	    RECT 2.3850 1.3450 2.6750 1.4000 ;
      END
   END SCE
   PIN SETB
      PORT
         LAYER li1 ;
	    RECT 6.5850 1.7850 7.0650 2.2950 ;
	    RECT 8.8800 1.9300 9.9450 2.1550 ;
	    RECT 8.8800 1.7800 9.1350 1.9300 ;
         LAYER met1 ;
	    RECT 6.5800 2.0000 6.8700 2.0550 ;
	    RECT 8.8800 2.0000 9.1700 2.0550 ;
	    RECT 6.5800 1.8250 9.1700 2.0000 ;
	    RECT 6.5800 1.7700 6.8700 1.8250 ;
	    RECT 8.8800 1.7700 9.1700 1.8250 ;
      END
   END SETB
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.1050 0.7000 0.7450 ;
	    RECT 1.8250 0.1050 2.0900 0.6800 ;
	    RECT 2.6900 0.1050 3.1000 0.6950 ;
	    RECT 3.6250 0.1050 3.9550 0.6800 ;
	    RECT 5.6100 0.1050 6.0950 0.5800 ;
	    RECT 6.7050 0.1050 7.7150 1.0050 ;
	    RECT 10.1150 0.1050 10.3650 0.6800 ;
	    RECT 11.5700 0.1050 11.8650 1.0300 ;
	    RECT 12.5350 0.1050 12.7950 1.1050 ;
	    RECT 0.0850 0.0850 12.7950 0.1050 ;
	    RECT 0.0000 -0.0850 12.8800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 12.8800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 12.8800 3.4850 ;
	    RECT 0.5150 3.2950 12.7950 3.3150 ;
	    RECT 0.5150 2.7450 0.7850 3.2950 ;
	    RECT 2.6900 2.6750 2.9850 3.2950 ;
	    RECT 3.5950 2.8450 3.9250 3.2950 ;
	    RECT 5.9450 2.8450 6.3300 3.2950 ;
	    RECT 7.0600 2.6550 8.0150 3.2950 ;
	    RECT 9.1600 2.7950 9.4900 3.2950 ;
	    RECT 10.1550 2.7950 10.4850 3.2950 ;
	    RECT 11.5700 2.2400 11.8200 3.2950 ;
	    RECT 12.5350 1.8700 12.7950 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 12.8800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.5300 0.3450 3.0800 ;
	    RECT 0.9550 2.8200 2.0450 3.0800 ;
	    RECT 0.9550 2.5300 1.1250 2.8200 ;
	    RECT 2.2700 2.6050 2.5200 3.0800 ;
	    RECT 0.0850 2.3050 1.1250 2.5300 ;
	    RECT 1.2950 2.3050 1.6950 2.6050 ;
	    RECT 1.5050 0.8900 1.6950 2.3050 ;
	    RECT 1.8650 2.2150 2.5200 2.6050 ;
	    RECT 3.2550 2.5000 3.4250 2.9050 ;
	    RECT 4.0950 2.6700 4.4400 3.0800 ;
	    RECT 3.2550 2.4900 3.9850 2.5000 ;
	    RECT 3.2550 2.2900 3.9950 2.4900 ;
	    RECT 1.8650 1.1300 2.2000 2.2150 ;
	    RECT 1.8650 0.8950 2.5200 1.1300 ;
	    RECT 3.7350 1.1050 3.9950 2.2900 ;
	    RECT 1.5050 0.8800 1.6750 0.8900 ;
	    RECT 1.4950 0.8300 1.6750 0.8800 ;
	    RECT 1.4750 0.8250 1.6750 0.8300 ;
	    RECT 1.4750 0.8050 1.6700 0.8250 ;
	    RECT 1.4600 0.7950 1.6650 0.8050 ;
	    RECT 1.4450 0.7900 1.6650 0.7950 ;
	    RECT 1.4400 0.7750 1.6650 0.7900 ;
	    RECT 1.4300 0.7700 1.6600 0.7750 ;
	    RECT 1.4200 0.7650 1.6600 0.7700 ;
	    RECT 1.4050 0.7550 1.6600 0.7650 ;
	    RECT 1.3950 0.7500 1.6600 0.7550 ;
	    RECT 1.3800 0.7450 1.6600 0.7500 ;
	    RECT 0.8700 0.7200 1.6500 0.7450 ;
	    RECT 0.8700 0.6950 1.6400 0.7200 ;
	    RECT 0.8700 0.3200 1.6250 0.6950 ;
	    RECT 2.2600 0.3200 2.5200 0.8950 ;
	    RECT 3.2700 0.8950 3.9950 1.1050 ;
	    RECT 4.1650 1.7750 4.4400 2.6700 ;
	    RECT 4.6150 2.0200 4.8300 3.0800 ;
	    RECT 5.0350 2.6700 5.7550 3.0800 ;
	    RECT 4.6150 1.9900 4.9150 2.0200 ;
	    RECT 4.6600 1.8050 4.9150 1.9900 ;
	    RECT 5.2050 1.9700 5.4150 2.4450 ;
	    RECT 4.1650 1.3650 4.4900 1.7750 ;
	    RECT 3.2700 0.3200 3.4550 0.8950 ;
	    RECT 4.1650 0.7300 4.3350 1.3650 ;
	    RECT 4.6600 1.1500 4.8300 1.8050 ;
	    RECT 5.5850 1.7450 5.7550 2.6700 ;
	    RECT 6.6050 2.6350 6.8200 3.0650 ;
	    RECT 8.1850 2.6550 8.9900 3.0750 ;
	    RECT 5.9250 2.4650 6.8200 2.6350 ;
	    RECT 8.8200 2.5800 8.9900 2.6550 ;
	    RECT 9.6600 2.5800 9.9650 3.0650 ;
	    RECT 5.9250 1.9700 6.0950 2.4650 ;
	    RECT 7.2350 2.0900 8.1350 2.4450 ;
	    RECT 5.0850 1.6550 5.7550 1.7450 ;
	    RECT 5.0850 1.6150 6.4750 1.6550 ;
	    RECT 7.3550 1.6150 7.7150 1.6550 ;
	    RECT 5.0850 1.5950 7.7150 1.6150 ;
	    RECT 4.1250 0.3200 4.3350 0.7300 ;
	    RECT 4.5050 0.3200 4.8300 1.1500 ;
	    RECT 5.0000 1.4450 7.7150 1.5950 ;
	    RECT 5.0000 0.3200 5.4400 1.4450 ;
	    RECT 5.6450 1.0050 5.9750 1.2700 ;
	    RECT 6.3050 1.2200 7.7150 1.4450 ;
	    RECT 7.8850 1.1300 8.1350 2.0900 ;
	    RECT 8.4250 1.3450 8.6500 2.3800 ;
	    RECT 8.8200 2.3700 10.4850 2.5800 ;
	    RECT 10.1550 2.0050 10.4850 2.3700 ;
	    RECT 10.6550 1.7050 10.9150 3.0800 ;
	    RECT 8.8200 1.1300 9.1050 1.5700 ;
	    RECT 5.6450 0.7950 6.5350 1.0050 ;
	    RECT 7.8850 0.9000 9.1050 1.1300 ;
	    RECT 9.3200 1.4950 10.9150 1.7050 ;
	    RECT 9.3200 1.0700 9.5300 1.4950 ;
	    RECT 9.7100 0.9800 10.5150 1.2700 ;
	    RECT 6.2850 0.3200 6.5350 0.7950 ;
	    RECT 9.7100 0.6800 9.9100 0.9800 ;
	    RECT 10.6850 0.7300 10.9150 1.4950 ;
	    RECT 8.4650 0.3450 9.9100 0.6800 ;
	    RECT 10.5750 0.3200 10.9150 0.7300 ;
	    RECT 11.0850 1.6550 11.3450 3.0800 ;
	    RECT 11.0850 1.2450 11.9750 1.6550 ;
	    RECT 11.0850 0.3200 11.3450 1.2450 ;
         LAYER met1 ;
	    RECT 3.7650 2.4250 4.0550 2.4800 ;
	    RECT 5.1450 2.4250 5.4350 2.4800 ;
	    RECT 7.5000 2.4250 7.7900 2.4800 ;
	    RECT 3.7650 2.2500 7.7900 2.4250 ;
	    RECT 3.7650 2.1950 4.0550 2.2500 ;
	    RECT 5.1450 2.1950 5.4350 2.2500 ;
	    RECT 7.5000 2.1950 7.7900 2.2500 ;
	    RECT 1.4650 2.0000 1.7550 2.0550 ;
	    RECT 4.6850 2.0000 4.9750 2.0550 ;
	    RECT 1.4650 1.8250 4.9750 2.0000 ;
	    RECT 1.4650 1.7700 1.7550 1.8250 ;
	    RECT 4.6850 1.7700 4.9750 1.8250 ;
	    RECT 4.2250 1.5750 4.5150 1.6300 ;
	    RECT 8.4200 1.5750 8.7100 1.6300 ;
	    RECT 4.2250 1.4000 8.7100 1.5750 ;
	    RECT 4.2250 1.3450 4.5150 1.4000 ;
	    RECT 8.4200 1.3450 8.7100 1.4000 ;
   END
END efs8hd_sdfstp_2
MACRO efs8hd_sdfxbp_2
   CLASS CORE ;
   FOREIGN efs8hd_sdfxbp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 11.9600 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.9750 0.1050 2.3050 0.5550 ;
	    RECT 3.7650 0.1050 3.9650 0.6550 ;
	    RECT 5.7150 0.1050 6.0850 0.7300 ;
	    RECT 7.7400 0.1050 8.1100 0.7700 ;
	    RECT 8.8950 0.1050 9.0850 0.8700 ;
	    RECT 9.7550 0.1050 9.9850 0.8650 ;
	    RECT 10.6900 0.1050 11.0200 1.0050 ;
	    RECT 11.6100 0.1050 11.7800 1.1950 ;
	    RECT 0.0000 -0.1050 11.9600 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 11.9600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 11.9600 3.5050 ;
	    RECT 0.5200 2.6700 0.8500 3.2950 ;
	    RECT 1.8800 2.8050 2.2100 3.2950 ;
	    RECT 3.7600 2.7050 3.9300 3.2950 ;
	    RECT 5.9250 2.2950 6.0950 3.2950 ;
	    RECT 7.8050 2.6700 8.1100 3.2950 ;
	    RECT 8.8950 2.0300 9.0750 3.2950 ;
	    RECT 9.7650 2.0200 9.9350 3.2950 ;
	    RECT 10.7150 1.8700 11.0200 3.2950 ;
	    RECT 11.6100 1.7450 11.7800 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 11.9600 3.7000 ;
      END
   END vpwr
   PIN SCD
      PORT
         LAYER li1 ;
	    RECT 3.5350 1.2950 4.0350 2.0700 ;
      END
   END SCD
   PIN D
      PORT
         LAYER li1 ;
	    RECT 2.4600 1.6950 2.7950 2.1050 ;
      END
   END D
   PIN QN
      PORT
         LAYER li1 ;
	    RECT 11.1900 1.8050 11.4400 2.9050 ;
	    RECT 11.2350 0.9950 11.4400 1.8050 ;
	    RECT 11.1900 0.3300 11.4400 0.9950 ;
      END
   END QN
   PIN SCE
      PORT
         LAYER li1 ;
	    RECT 1.7800 0.9800 1.9500 2.1050 ;
	    RECT 3.0850 0.9800 3.2550 1.3950 ;
	    RECT 1.7800 0.7700 3.2550 0.9800 ;
	    RECT 2.4750 0.3800 2.6500 0.7700 ;
      END
   END SCE
   PIN CLK
      PORT
         LAYER li1 ;
	    RECT 0.0950 1.2200 0.4450 2.0300 ;
      END
   END CLK
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 9.2550 1.9150 9.5850 3.0400 ;
	    RECT 9.2550 1.8700 9.6150 1.9150 ;
	    RECT 9.4100 1.7900 9.6150 1.8700 ;
	    RECT 9.4450 1.1150 9.6150 1.7900 ;
	    RECT 9.4100 1.0300 9.6150 1.1150 ;
	    RECT 9.2550 0.9900 9.6150 1.0300 ;
	    RECT 9.2550 0.3200 9.5850 0.9900 ;
      END
   END Q
   OBS
         LAYER li1 ;
	    RECT 0.1800 2.4550 0.3500 3.0800 ;
	    RECT 0.1800 2.2450 0.8450 2.4550 ;
	    RECT 0.6150 1.2150 0.8450 2.2450 ;
	    RECT 0.6150 1.0050 0.8100 1.2150 ;
	    RECT 0.1750 0.7950 0.8100 1.0050 ;
	    RECT 1.0200 0.8950 1.2450 3.0800 ;
	    RECT 0.1750 0.4300 0.3450 0.7950 ;
	    RECT 1.0150 0.4300 1.2450 0.8950 ;
	    RECT 1.4350 2.5950 1.7100 3.0550 ;
	    RECT 2.6950 2.8050 3.5900 3.0200 ;
	    RECT 1.4350 2.3250 3.2500 2.5950 ;
	    RECT 1.4350 0.5550 1.6050 2.3250 ;
	    RECT 2.1200 1.4050 2.2900 2.3250 ;
	    RECT 3.0800 2.1050 3.2500 2.3250 ;
	    RECT 3.4200 2.4950 3.5900 2.8050 ;
	    RECT 4.2050 2.5800 4.4850 3.0500 ;
	    RECT 4.6850 2.7400 5.7550 2.9500 ;
	    RECT 4.2050 2.4950 4.3750 2.5800 ;
	    RECT 3.4200 2.2800 4.3750 2.4950 ;
	    RECT 3.0800 1.6950 3.2750 2.1050 ;
	    RECT 2.1200 1.1950 2.4650 1.4050 ;
	    RECT 4.2050 1.0800 4.3750 2.2800 ;
	    RECT 3.4250 0.8700 4.3750 1.0800 ;
	    RECT 4.5450 1.2950 4.7850 2.3800 ;
	    RECT 4.9750 2.0700 5.4150 2.5150 ;
	    RECT 5.5850 1.9700 5.7550 2.7400 ;
	    RECT 6.2650 2.6700 6.5150 3.0800 ;
	    RECT 6.7400 2.7050 7.6250 2.9200 ;
	    RECT 5.5850 1.8550 6.0950 1.9700 ;
	    RECT 5.2950 1.6450 6.0950 1.8550 ;
	    RECT 4.5450 0.8800 5.1250 1.2950 ;
	    RECT 3.4250 0.5550 3.5950 0.8700 ;
	    RECT 1.4350 0.3450 1.8050 0.5550 ;
	    RECT 2.8200 0.3450 3.5950 0.5550 ;
	    RECT 4.2050 0.6700 4.3750 0.8700 ;
	    RECT 5.2950 0.6700 5.4650 1.6450 ;
	    RECT 5.9250 1.5550 6.0950 1.6450 ;
	    RECT 5.6350 1.3300 5.8050 1.3700 ;
	    RECT 6.2650 1.3300 6.4350 2.6700 ;
	    RECT 6.6050 1.5550 6.7950 2.4550 ;
	    RECT 6.9650 1.9700 7.2850 2.3800 ;
	    RECT 5.6350 0.9550 6.4350 1.3300 ;
	    RECT 6.9650 1.2950 7.1550 1.9700 ;
	    RECT 7.4550 1.7550 7.6250 2.7050 ;
	    RECT 8.3950 2.3800 8.7250 3.0700 ;
	    RECT 7.7950 1.9700 8.7250 2.3800 ;
	    RECT 4.2050 0.4550 4.5550 0.6700 ;
	    RECT 4.7250 0.4550 5.4650 0.6700 ;
	    RECT 6.2650 0.6700 6.4350 0.9550 ;
	    RECT 6.6050 0.8800 7.1550 1.2950 ;
	    RECT 7.3250 1.6550 7.6250 1.7550 ;
	    RECT 8.5400 1.6550 8.7250 1.9700 ;
	    RECT 10.2050 1.6550 10.5350 3.0300 ;
	    RECT 7.3250 1.2450 8.3700 1.6550 ;
	    RECT 8.5400 1.2450 9.2750 1.6550 ;
	    RECT 10.2050 1.2450 11.0650 1.6550 ;
	    RECT 7.3250 0.6700 7.4950 1.2450 ;
	    RECT 8.5400 1.0300 8.7250 1.2450 ;
	    RECT 6.2650 0.4550 6.7250 0.6700 ;
	    RECT 6.9550 0.4550 7.4950 0.6700 ;
	    RECT 8.3600 0.3750 8.7250 1.0300 ;
	    RECT 10.2050 0.4300 10.4550 1.2450 ;
         LAYER met1 ;
	    RECT 0.5850 2.4250 0.8750 2.4800 ;
	    RECT 5.1450 2.4250 5.4350 2.4800 ;
	    RECT 6.5650 2.4250 6.8550 2.4800 ;
	    RECT 0.5850 2.2500 6.8550 2.4250 ;
	    RECT 0.5850 2.1950 0.8750 2.2500 ;
	    RECT 5.1450 2.1950 5.4350 2.2500 ;
	    RECT 6.5650 2.1950 6.8550 2.2500 ;
	    RECT 0.9900 1.1500 1.2800 1.2050 ;
	    RECT 4.6850 1.1500 4.9750 1.2050 ;
	    RECT 6.5800 1.1500 6.8700 1.2050 ;
	    RECT 0.9900 0.9750 6.8700 1.1500 ;
	    RECT 0.9900 0.9200 1.2800 0.9750 ;
	    RECT 4.6850 0.9200 4.9750 0.9750 ;
	    RECT 6.5800 0.9200 6.8700 0.9750 ;
   END
END efs8hd_sdfxbp_2
MACRO efs8hd_sdfxtp_2
   CLASS CORE ;
   FOREIGN efs8hd_sdfxtp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 10.1200 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5800 ;
	    RECT 1.9750 0.1050 2.3050 0.5550 ;
	    RECT 3.7600 0.1050 3.9600 0.6550 ;
	    RECT 5.7200 0.1050 6.0900 0.7300 ;
	    RECT 7.7450 0.1050 8.1150 0.7700 ;
	    RECT 8.9050 0.1050 9.0750 0.8700 ;
	    RECT 9.7750 0.1050 9.9450 1.1650 ;
	    RECT 0.0000 -0.1050 10.1200 0.1050 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 10.1200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.2950 10.1200 3.5050 ;
	    RECT 0.5200 2.6700 0.8500 3.2950 ;
	    RECT 1.8800 2.8050 2.2100 3.2950 ;
	    RECT 3.7550 2.7050 3.9250 3.2950 ;
	    RECT 5.9300 2.2950 6.1000 3.2950 ;
	    RECT 7.8100 2.6700 8.1150 3.2950 ;
	    RECT 8.9050 2.0300 9.0800 3.2950 ;
	    RECT 9.7750 1.7550 9.9450 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 10.1200 3.7000 ;
      END
   END vpwr
   PIN SCD
      PORT
         LAYER li1 ;
	    RECT 3.5300 1.2950 4.0200 2.0700 ;
      END
   END SCD
   PIN D
      PORT
         LAYER li1 ;
	    RECT 2.4600 1.6950 2.7900 2.1050 ;
      END
   END D
   PIN SCE
      PORT
         LAYER li1 ;
	    RECT 1.7800 0.9800 1.9500 2.1050 ;
	    RECT 3.0800 0.9800 3.2500 1.3950 ;
	    RECT 1.7800 0.7700 3.2500 0.9800 ;
	    RECT 2.4750 0.3800 2.6500 0.7700 ;
      END
   END SCE
   PIN CLK
      PORT
         LAYER li1 ;
	    RECT 0.0950 1.2200 0.4450 2.0300 ;
      END
   END CLK
   PIN Q
      PORT
         LAYER li1 ;
	    RECT 9.2600 1.8800 9.6050 2.9950 ;
	    RECT 9.4350 1.0250 9.6050 1.8800 ;
	    RECT 9.2600 0.3800 9.6050 1.0250 ;
      END
   END Q
   OBS
         LAYER li1 ;
	    RECT 0.1800 2.4550 0.3500 3.0800 ;
	    RECT 0.1800 2.2450 0.8450 2.4550 ;
	    RECT 0.6150 1.2150 0.8450 2.2450 ;
	    RECT 0.6150 1.0050 0.8100 1.2150 ;
	    RECT 0.1750 0.7950 0.8100 1.0050 ;
	    RECT 1.0200 0.8950 1.2450 3.0800 ;
	    RECT 0.1750 0.4300 0.3450 0.7950 ;
	    RECT 1.0150 0.4300 1.2450 0.8950 ;
	    RECT 1.4350 2.5950 1.7100 3.0550 ;
	    RECT 2.6900 2.8050 3.5850 3.0200 ;
	    RECT 1.4350 2.3250 3.2450 2.5950 ;
	    RECT 1.4350 0.5550 1.6050 2.3250 ;
	    RECT 2.1200 1.4050 2.2900 2.3250 ;
	    RECT 3.0750 2.1050 3.2450 2.3250 ;
	    RECT 3.4150 2.4950 3.5850 2.8050 ;
	    RECT 4.2100 2.5800 4.4450 3.0500 ;
	    RECT 4.6900 2.7400 5.7600 2.9500 ;
	    RECT 4.2100 2.4950 4.3800 2.5800 ;
	    RECT 3.4150 2.2800 4.3800 2.4950 ;
	    RECT 3.0750 1.6950 3.2700 2.1050 ;
	    RECT 2.1200 1.1950 2.4600 1.4050 ;
	    RECT 4.2100 1.0800 4.3800 2.2800 ;
	    RECT 3.4200 0.8700 4.3800 1.0800 ;
	    RECT 4.5500 1.2950 4.7900 2.3800 ;
	    RECT 4.9800 2.0700 5.4200 2.5150 ;
	    RECT 5.5900 1.9700 5.7600 2.7400 ;
	    RECT 6.2700 2.6700 6.5200 3.0800 ;
	    RECT 6.7450 2.7050 7.6300 2.9200 ;
	    RECT 5.5900 1.8550 6.1000 1.9700 ;
	    RECT 5.3000 1.6450 6.1000 1.8550 ;
	    RECT 4.5500 0.8800 5.1300 1.2950 ;
	    RECT 3.4200 0.5550 3.5900 0.8700 ;
	    RECT 1.4350 0.3450 1.8050 0.5550 ;
	    RECT 2.8200 0.3450 3.5900 0.5550 ;
	    RECT 4.2100 0.6700 4.3800 0.8700 ;
	    RECT 5.3000 0.6700 5.4700 1.6450 ;
	    RECT 5.9300 1.5550 6.1000 1.6450 ;
	    RECT 5.6400 1.3300 5.8100 1.3700 ;
	    RECT 6.2700 1.3300 6.4400 2.6700 ;
	    RECT 6.6100 1.5550 6.8000 2.4550 ;
	    RECT 6.9700 1.9700 7.2900 2.3800 ;
	    RECT 5.6400 0.9550 6.4400 1.3300 ;
	    RECT 6.9700 1.2950 7.1600 1.9700 ;
	    RECT 7.4600 1.7550 7.6300 2.7050 ;
	    RECT 8.4650 2.3800 8.7350 3.0700 ;
	    RECT 7.8000 1.9700 8.7350 2.3800 ;
	    RECT 4.2100 0.4550 4.5600 0.6700 ;
	    RECT 4.7300 0.4550 5.4700 0.6700 ;
	    RECT 6.2700 0.6700 6.4400 0.9550 ;
	    RECT 6.6100 0.8800 7.1600 1.2950 ;
	    RECT 7.3300 1.6550 7.6300 1.7550 ;
	    RECT 8.5650 1.6550 8.7350 1.9700 ;
	    RECT 7.3300 1.2450 8.3950 1.6550 ;
	    RECT 8.5650 1.2450 9.2650 1.6550 ;
	    RECT 7.3300 0.6700 7.5000 1.2450 ;
	    RECT 8.5650 1.0300 8.7350 1.2450 ;
	    RECT 6.2700 0.4550 6.7300 0.6700 ;
	    RECT 6.9600 0.4550 7.5000 0.6700 ;
	    RECT 8.3850 0.3750 8.7350 1.0300 ;
         LAYER met1 ;
	    RECT 0.5800 2.4250 0.8700 2.4800 ;
	    RECT 5.1450 2.4250 5.4350 2.4800 ;
	    RECT 6.5600 2.4250 6.8500 2.4800 ;
	    RECT 0.5800 2.2500 6.8500 2.4250 ;
	    RECT 0.5800 2.1950 0.8700 2.2500 ;
	    RECT 5.1450 2.1950 5.4350 2.2500 ;
	    RECT 6.5600 2.1950 6.8500 2.2500 ;
	    RECT 0.9900 1.1500 1.2800 1.2050 ;
	    RECT 4.6850 1.1500 4.9750 1.2050 ;
	    RECT 6.5700 1.1500 6.8600 1.2050 ;
	    RECT 0.9900 0.9750 6.8600 1.1500 ;
	    RECT 0.9900 0.9200 1.2800 0.9750 ;
	    RECT 4.6850 0.9200 4.9750 0.9750 ;
	    RECT 6.5700 0.9200 6.8600 0.9750 ;
   END
END efs8hd_sdfxtp_2
MACRO efs8hd_sdlclkp_2
   CLASS CORE ;
   FOREIGN efs8hd_sdlclkp_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 7.3600 BY 3.4000 ;
   SITE unitehd ;
   PIN GCLK
      PORT
         LAYER li1 ;
	    RECT 6.5700 1.8700 6.8400 3.0800 ;
	    RECT 6.6700 1.6450 6.8400 1.8700 ;
	    RECT 6.6700 1.3200 7.2750 1.6450 ;
	    RECT 6.6700 1.0300 6.8400 1.3200 ;
	    RECT 6.5700 0.3200 6.8400 1.0300 ;
      END
   END GCLK
   PIN SCE
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.1050 0.3400 2.0800 ;
      END
   END SCE
   PIN CLK
      PORT
         LAYER li1 ;
	    RECT 4.7050 1.6150 4.9250 1.6550 ;
	    RECT 4.7050 1.1950 6.0500 1.6150 ;
      END
   END CLK
   PIN GATE
      PORT
         LAYER li1 ;
	    RECT 0.8550 1.8050 1.2400 2.4450 ;
	    RECT 0.8550 1.1950 1.2350 1.8050 ;
      END
   END GATE
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.8450 0.5550 ;
	    RECT 2.6700 0.1050 3.0150 1.0300 ;
	    RECT 4.0950 0.1050 4.4250 0.5550 ;
	    RECT 5.4900 0.1050 6.4000 0.5550 ;
	    RECT 7.0100 0.1050 7.2750 1.1050 ;
	    RECT 0.5150 0.0850 7.2750 0.1050 ;
	    RECT 0.0000 -0.0850 7.3600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 7.3600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 7.3600 3.4850 ;
	    RECT 0.0850 3.2950 7.2750 3.3150 ;
	    RECT 0.0850 2.2950 0.3450 3.2950 ;
	    RECT 2.3750 2.5950 3.0150 3.2950 ;
	    RECT 3.5750 2.8200 5.5300 3.2950 ;
	    RECT 6.0700 2.8200 6.4000 3.2950 ;
	    RECT 7.0100 1.8550 7.2750 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 7.3600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.5150 2.6550 1.2600 3.0800 ;
	    RECT 1.4300 2.6550 2.2050 3.0800 ;
	    RECT 0.5150 0.9800 0.6850 2.6550 ;
	    RECT 1.4100 1.6550 1.8650 2.4450 ;
	    RECT 1.4050 1.5050 1.8650 1.6550 ;
	    RECT 2.0350 1.7200 2.2050 2.6550 ;
	    RECT 3.1850 2.6050 3.4050 3.0800 ;
	    RECT 5.7000 2.6050 5.8700 3.0800 ;
	    RECT 3.1850 2.3950 5.4900 2.6050 ;
	    RECT 3.1850 2.3800 3.4050 2.3950 ;
	    RECT 2.3750 2.0450 3.4050 2.3800 ;
	    RECT 2.3750 1.9700 2.5450 2.0450 ;
	    RECT 2.0350 1.5050 3.0150 1.7200 ;
	    RECT 0.5150 0.9350 1.1950 0.9800 ;
	    RECT 0.0850 0.7650 1.1950 0.9350 ;
	    RECT 1.4050 0.8800 1.7050 1.5050 ;
	    RECT 1.8750 0.8800 2.1600 1.2950 ;
	    RECT 2.3300 1.2450 3.0150 1.5050 ;
	    RECT 0.0850 0.3200 0.3450 0.7650 ;
	    RECT 1.0150 0.3200 1.1950 0.7650 ;
	    RECT 2.3300 0.6700 2.5000 1.2450 ;
	    RECT 1.3650 0.3200 2.5000 0.6700 ;
	    RECT 3.1850 0.3200 3.4050 2.0450 ;
	    RECT 3.5750 1.9700 4.0400 2.1800 ;
	    RECT 3.5750 1.1700 3.7450 1.9700 ;
	    RECT 4.2100 1.8700 5.0100 2.1800 ;
	    RECT 5.1800 2.0050 5.4900 2.3950 ;
	    RECT 5.7000 2.2200 6.4000 2.6050 ;
	    RECT 4.2100 1.5950 4.4600 1.8700 ;
	    RECT 5.1800 1.7950 5.6500 2.0050 ;
	    RECT 5.8200 1.7950 6.4000 2.2200 ;
	    RECT 3.9150 1.3800 4.4600 1.5950 ;
	    RECT 3.5750 0.9550 4.0000 1.1700 ;
	    RECT 4.1700 0.9800 4.4600 1.3800 ;
	    RECT 6.2300 1.6550 6.4000 1.7950 ;
	    RECT 6.2300 1.2450 6.5000 1.6550 ;
	    RECT 6.2300 0.9800 6.4000 1.2450 ;
	    RECT 3.5750 0.3200 3.9250 0.9550 ;
	    RECT 4.1700 0.7700 4.8250 0.9800 ;
	    RECT 4.5950 0.3200 4.8250 0.7700 ;
	    RECT 5.1000 0.7700 6.4000 0.9800 ;
	    RECT 5.1000 0.3200 5.3100 0.7700 ;
         LAYER met1 ;
	    RECT 1.4700 2.0000 1.7600 2.0550 ;
	    RECT 4.2300 2.0000 4.5200 2.0550 ;
	    RECT 1.4700 1.8250 4.5200 2.0000 ;
	    RECT 1.4700 1.7700 1.7600 1.8250 ;
	    RECT 4.2300 1.7700 4.5200 1.8250 ;
	    RECT 1.9300 1.1500 2.2200 1.2050 ;
	    RECT 3.7700 1.1500 4.0600 1.2050 ;
	    RECT 1.9300 0.9750 4.0600 1.1500 ;
	    RECT 1.9300 0.9200 2.2200 0.9750 ;
	    RECT 3.7700 0.9200 4.0600 0.9750 ;
   END
END efs8hd_sdlclkp_2
MACRO efs8hd_tap_1
   CLASS CORE ;
   FOREIGN efs8hd_tap_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 0.4600 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0000 -0.0850 0.4600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 0.4600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 0.4600 3.4850 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 0.4600 3.7000 ;
      END
   END vpwr
   PIN vnb
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.3300 0.3750 1.0100 ;
      END
   END vnb
   PIN vpb
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.8350 0.3750 3.0650 ;
      END
   END vpb
END efs8hd_tap_1
MACRO efs8hd_tap_2
   CLASS CORE ;
   FOREIGN efs8hd_tap_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 0.9200 BY 3.4000 ;
   SITE unitehd ;
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0000 -0.0850 0.9200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 0.9200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 0.9200 3.4850 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 0.9200 3.7000 ;
      END
   END vpwr
   PIN vpb
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.8350 0.8350 3.0650 ;
      END
   END vpb
   PIN vnb
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.3300 0.8350 1.0100 ;
      END
   END vnb
END efs8hd_tap_2
MACRO efs8hd_tapvgnd_1
   CLASS CORE ;
   FOREIGN efs8hd_tapvgnd_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 0.4600 BY 3.4000 ;
   SITE unitehd ;
   PIN vpb
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.8350 0.3750 3.0650 ;
         LAYER met1 ;
	    RECT 0.0850 2.6150 0.3750 2.9050 ;
      END
   END vpb
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.0850 0.3750 1.0100 ;
	    RECT 0.0000 -0.0850 0.4600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 0.4600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 0.4600 3.4850 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 0.4600 3.7000 ;
      END
   END vpwr
END efs8hd_tapvgnd_1
MACRO efs8hd_tapvgnd2_1
   CLASS CORE ;
   FOREIGN efs8hd_tapvgnd2_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 0.4600 BY 3.4000 ;
   SITE unitehd ;
   PIN vpb
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.8350 0.3750 3.0650 ;
         LAYER met1 ;
	    RECT 0.0850 2.1900 0.3750 2.4800 ;
      END
   END vpb
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.0850 0.3750 1.0100 ;
	    RECT 0.0000 -0.0850 0.4600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 0.4600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 0.4600 3.4850 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 0.4600 3.7000 ;
      END
   END vpwr
END efs8hd_tapvgnd2_1
MACRO efs8hd_tapvpwrvgnd_1
   CLASS CORE ;
   FOREIGN efs8hd_tapvpwrvgnd_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 0.4600 BY 3.4000 ;
   SITE unitehd ;
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 0.4600 3.4850 ;
	    RECT 0.0850 1.8350 0.3750 3.3150 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 0.4600 3.7000 ;
      END
   END vpwr
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.0850 0.3750 1.0100 ;
	    RECT 0.0000 -0.0850 0.4600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 0.4600 0.3000 ;
      END
   END vgnd
END efs8hd_tapvpwrvgnd_1
MACRO efs8hd_xnor2_2
   CLASS CORE ;
   FOREIGN efs8hd_xnor2_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.9800 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 1.2550 1.3450 2.7050 1.6150 ;
      END
   END A
   PIN B
      PORT
         LAYER li1 ;
	    RECT 0.7900 1.7850 3.1000 2.0200 ;
	    RECT 0.7900 1.6050 0.9600 1.7850 ;
	    RECT 0.4850 1.3450 0.9600 1.6050 ;
	    RECT 2.9300 1.6050 3.1000 1.7850 ;
	    RECT 2.9300 1.3450 3.9550 1.6050 ;
      END
   END B
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 3.7250 2.4550 3.9350 2.6550 ;
	    RECT 5.0450 2.4550 5.2950 2.6550 ;
	    RECT 3.7250 2.2450 5.2950 2.4550 ;
	    RECT 5.0450 2.0300 5.2950 2.2450 ;
	    RECT 5.0450 1.7700 5.8950 2.0300 ;
	    RECT 5.5050 0.5950 5.8950 1.7700 ;
	    RECT 4.5850 0.3800 5.8950 0.5950 ;
      END
   END Y
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 1.4500 0.1050 1.6200 0.6950 ;
	    RECT 2.4300 0.1050 2.6000 1.1300 ;
	    RECT 3.2700 0.1050 3.4400 0.6950 ;
	    RECT 4.1450 0.1050 4.3150 0.6950 ;
	    RECT 1.4500 0.0850 4.3150 0.1050 ;
	    RECT 0.0000 -0.0850 5.9800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.9800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.9800 3.4850 ;
	    RECT 0.5700 3.2950 5.8950 3.3150 ;
	    RECT 0.5700 2.6700 0.8200 3.2950 ;
	    RECT 1.4100 2.6700 1.6600 3.2950 ;
	    RECT 2.8100 2.6700 3.0600 3.2950 ;
	    RECT 4.6250 2.6700 4.8750 3.2950 ;
	    RECT 5.4650 2.2450 5.8950 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.9800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.4550 0.4000 3.0800 ;
	    RECT 0.9900 2.4550 1.2400 3.0800 ;
	    RECT 1.8300 2.4550 2.0800 3.0800 ;
	    RECT 2.3900 2.6550 2.6400 3.0800 ;
	    RECT 3.2300 2.8700 4.3550 3.0800 ;
	    RECT 3.2300 2.6550 3.5550 2.8700 ;
	    RECT 4.1050 2.6700 4.3550 2.8700 ;
	    RECT 0.0850 2.4450 2.0800 2.4550 ;
	    RECT 0.0850 2.2300 3.4800 2.4450 ;
	    RECT 0.0850 1.1200 0.3150 2.2300 ;
	    RECT 3.3100 2.0300 3.4800 2.2300 ;
	    RECT 3.3100 1.8200 4.8050 2.0300 ;
	    RECT 4.6350 1.5550 4.8050 1.8200 ;
	    RECT 4.6350 1.3450 5.2950 1.5550 ;
	    RECT 0.0850 0.8050 0.8600 1.1200 ;
	    RECT 1.0300 0.9050 2.1200 1.1300 ;
	    RECT 1.0300 0.5950 1.2800 0.9050 ;
	    RECT 0.1050 0.3200 1.2800 0.5950 ;
	    RECT 1.7900 0.3200 2.1200 0.9050 ;
	    RECT 2.7700 0.9050 5.3350 1.1300 ;
	    RECT 2.7700 0.3200 3.1000 0.9050 ;
	    RECT 3.6100 0.3200 3.9750 0.9050 ;
	    RECT 5.0050 0.8050 5.3350 0.9050 ;
         LAYER met1 ;
	    RECT 2.4050 2.8500 2.6950 2.9050 ;
	    RECT 3.3250 2.8500 3.6150 2.9050 ;
	    RECT 2.4050 2.6750 3.6150 2.8500 ;
	    RECT 2.4050 2.6200 2.6950 2.6750 ;
	    RECT 3.3250 2.6200 3.6150 2.6750 ;
   END
END efs8hd_xnor2_2
MACRO efs8hd_xnor2_4
   CLASS CORE ;
   FOREIGN efs8hd_xnor2_4 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 10.1200 BY 3.4000 ;
   SITE unitehd ;
   PIN B
      PORT
         LAYER li1 ;
	    RECT 1.6850 1.7850 5.7300 2.0200 ;
	    RECT 1.6850 1.5950 1.8550 1.7850 ;
	    RECT 0.4900 1.3450 1.8550 1.5950 ;
	    RECT 5.5600 1.5950 5.7300 1.7850 ;
	    RECT 5.5600 1.3450 7.4300 1.5950 ;
      END
   END B
   PIN A
      PORT
         LAYER li1 ;
	    RECT 2.1750 1.3450 5.3900 1.6150 ;
      END
   END A
   PIN Y
      PORT
         LAYER li1 ;
	    RECT 7.9600 2.5550 8.2500 3.0800 ;
	    RECT 6.1600 2.2300 8.2500 2.5550 ;
	    RECT 7.9600 2.0800 8.2500 2.2300 ;
	    RECT 8.8400 2.0800 9.0900 3.0800 ;
	    RECT 9.6800 2.0800 10.0350 3.0800 ;
	    RECT 7.9600 1.8050 10.0350 2.0800 ;
	    RECT 9.8150 1.1300 10.0350 1.8050 ;
	    RECT 8.3800 0.8050 10.0350 1.1300 ;
      END
   END Y
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 2.3500 0.1050 2.5200 0.6950 ;
	    RECT 3.1900 0.1050 3.3600 0.6950 ;
	    RECT 4.0350 0.1050 4.3100 1.1300 ;
	    RECT 4.9800 0.1050 5.1500 0.6950 ;
	    RECT 5.8200 0.1050 5.9900 0.6950 ;
	    RECT 6.6600 0.1050 6.8300 0.6950 ;
	    RECT 7.5000 0.1050 7.7700 0.6950 ;
	    RECT 2.3500 0.0850 7.7700 0.1050 ;
	    RECT 0.0000 -0.0850 10.1200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 10.1200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 10.1200 3.4850 ;
	    RECT 0.6300 3.2950 9.5100 3.3150 ;
	    RECT 0.6300 2.2950 0.8800 3.2950 ;
	    RECT 1.4700 2.7200 1.7200 3.2950 ;
	    RECT 2.3100 2.7200 2.5600 3.2950 ;
	    RECT 3.1500 2.7200 3.4000 3.2950 ;
	    RECT 4.5200 2.7200 4.7700 3.2950 ;
	    RECT 5.3600 2.7200 5.6100 3.2950 ;
	    RECT 8.4200 2.2950 8.6700 3.2950 ;
	    RECT 9.2600 2.2950 9.5100 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 10.1200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.0200 0.4600 3.0800 ;
	    RECT 1.0500 2.5050 1.3000 3.0800 ;
	    RECT 1.8900 2.5050 2.1400 3.0800 ;
	    RECT 2.7300 2.5050 2.9800 3.0800 ;
	    RECT 3.5700 2.5050 3.8200 3.0800 ;
	    RECT 1.0500 2.2300 3.8200 2.5050 ;
	    RECT 4.0350 2.5050 4.3500 3.0800 ;
	    RECT 4.9400 2.5050 5.1900 3.0800 ;
	    RECT 5.7800 2.7700 7.7500 3.0800 ;
	    RECT 5.7800 2.5050 5.9900 2.7700 ;
	    RECT 4.0350 2.2300 5.9900 2.5050 ;
	    RECT 1.0500 2.0200 1.3000 2.2300 ;
	    RECT 0.0850 1.8050 1.3000 2.0200 ;
	    RECT 5.9000 1.8050 7.7700 2.0200 ;
	    RECT 0.0850 1.1300 0.3200 1.8050 ;
	    RECT 7.6000 1.5950 7.7700 1.8050 ;
	    RECT 7.6000 1.3450 9.6450 1.5950 ;
	    RECT 0.0850 0.8050 1.7600 1.1300 ;
	    RECT 1.9300 0.9050 3.8600 1.1300 ;
	    RECT 1.9300 0.5950 2.1800 0.9050 ;
	    RECT 0.1700 0.3200 2.1800 0.5950 ;
	    RECT 2.6900 0.3200 3.0200 0.9050 ;
	    RECT 3.5300 0.3200 3.8600 0.9050 ;
	    RECT 4.4800 0.9200 8.2100 1.1300 ;
	    RECT 4.4800 0.9050 7.4300 0.9200 ;
	    RECT 4.4800 0.3200 4.8100 0.9050 ;
	    RECT 5.3200 0.3200 5.6500 0.9050 ;
	    RECT 6.1600 0.3200 6.4900 0.9050 ;
	    RECT 7.0000 0.3200 7.3300 0.9050 ;
	    RECT 7.9600 0.5950 8.2100 0.9200 ;
	    RECT 7.9600 0.3800 9.9700 0.5950 ;
         LAYER met1 ;
	    RECT 1.0050 2.0000 1.2950 2.0550 ;
	    RECT 6.0650 2.0000 6.3550 2.0550 ;
	    RECT 1.0050 1.8250 6.3550 2.0000 ;
	    RECT 1.0050 1.7700 1.2950 1.8250 ;
	    RECT 6.0650 1.7700 6.3550 1.8250 ;
   END
END efs8hd_xnor2_4
MACRO efs8hd_xnor3_1
   CLASS CORE ;
   FOREIGN efs8hd_xnor3_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 8.2800 BY 3.4000 ;
   SITE unitehd ;
   PIN C
      PORT
         LAYER li1 ;
	    RECT 1.6150 1.3450 2.1800 1.6550 ;
      END
   END C
   PIN A
      PORT
         LAYER li1 ;
	    RECT 7.0450 1.3450 7.4550 1.6550 ;
      END
   END A
   PIN B
      PORT
         LAYER li1 ;
	    RECT 6.1250 1.7850 6.8050 2.0200 ;
	    RECT 6.1250 1.2450 6.3950 1.7850 ;
      END
   END B
   PIN X
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.8000 0.3650 3.0800 ;
	    RECT 0.0850 1.1550 0.3300 1.8000 ;
	    RECT 0.0850 0.4400 0.3450 1.1550 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5150 0.1050 0.7650 0.6550 ;
	    RECT 3.4750 0.1050 3.6450 1.0800 ;
	    RECT 7.4750 0.1050 7.6450 0.7050 ;
	    RECT 0.5150 0.0850 7.6450 0.1050 ;
	    RECT 0.0000 -0.0850 8.2800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 8.2800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 8.2800 3.4850 ;
	    RECT 0.5350 3.2950 7.7300 3.3150 ;
	    RECT 0.5350 2.7700 0.8700 3.2950 ;
	    RECT 3.2250 2.7950 3.5550 3.2950 ;
	    RECT 7.3950 2.8450 7.7300 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 8.2800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 1.0500 2.7950 2.5200 3.0050 ;
	    RECT 3.8900 2.8450 6.9850 3.0550 ;
	    RECT 1.0500 2.5550 1.2200 2.7950 ;
	    RECT 3.8900 2.5800 4.0600 2.8450 ;
	    RECT 0.5350 2.3450 1.2200 2.5550 ;
	    RECT 1.5600 2.3700 4.0600 2.5800 ;
	    RECT 0.5350 1.6550 0.7050 2.3450 ;
	    RECT 0.9350 1.9200 2.5200 2.1300 ;
	    RECT 0.5000 1.2450 0.7050 1.6550 ;
	    RECT 0.5300 1.0800 0.7050 1.2450 ;
	    RECT 0.5300 0.8700 1.1050 1.0800 ;
	    RECT 0.9350 0.5300 1.1050 0.8700 ;
	    RECT 1.2750 0.7450 1.4450 1.9200 ;
	    RECT 2.3500 1.6550 2.5200 1.9200 ;
	    RECT 2.6900 1.9050 3.0750 2.1200 ;
	    RECT 2.7950 1.7200 3.0750 1.9050 ;
	    RECT 2.3500 1.2450 2.6250 1.6550 ;
	    RECT 1.7450 0.9950 2.1250 1.1300 ;
	    RECT 2.7950 0.9950 2.9650 1.7200 ;
	    RECT 3.2450 1.5050 3.4150 2.3700 ;
	    RECT 3.6450 1.8050 4.0650 2.1450 ;
	    RECT 1.7450 0.7800 2.9650 0.9950 ;
	    RECT 3.1350 1.2950 3.4150 1.5050 ;
	    RECT 3.1350 0.5700 3.3050 1.2950 ;
	    RECT 2.0700 0.5300 2.5050 0.5700 ;
	    RECT 0.9350 0.3200 2.5050 0.5300 ;
	    RECT 2.6750 0.3550 3.3050 0.5700 ;
	    RECT 3.8250 0.5200 4.0650 1.8050 ;
	    RECT 4.2450 0.7450 4.4150 2.6300 ;
	    RECT 4.5850 1.0750 4.7550 2.8450 ;
	    RECT 7.9000 2.6300 8.1950 3.0800 ;
	    RECT 4.9350 2.0200 5.3500 2.5550 ;
	    RECT 5.7850 2.4200 8.1950 2.6300 ;
	    RECT 4.9350 1.8050 5.6150 2.0200 ;
	    RECT 4.9500 1.2450 5.2750 1.5950 ;
	    RECT 4.5850 0.9000 4.9350 1.0750 ;
	    RECT 5.1050 0.9900 5.2750 1.2450 ;
	    RECT 4.6250 0.8550 4.9350 0.9000 ;
	    RECT 4.2450 0.5550 4.4550 0.7450 ;
	    RECT 4.6250 0.7250 4.9950 0.8550 ;
	    RECT 4.2450 0.3300 4.6550 0.5550 ;
	    RECT 4.8250 0.4000 4.9950 0.7250 ;
	    RECT 5.4450 0.5300 5.6150 1.8050 ;
	    RECT 5.7850 0.7450 5.9550 2.4200 ;
	    RECT 7.7100 2.3450 8.1950 2.4200 ;
	    RECT 6.9750 1.8700 7.7950 2.1300 ;
	    RECT 7.6250 1.6550 7.7950 1.8700 ;
	    RECT 6.5650 1.1800 6.8750 1.5950 ;
	    RECT 7.6250 1.2450 7.8550 1.6550 ;
	    RECT 6.5650 0.9150 6.7700 1.1800 ;
	    RECT 7.6250 1.1300 7.7950 1.2450 ;
	    RECT 7.0550 0.9400 7.7950 1.1300 ;
	    RECT 7.0150 0.9200 7.7950 0.9400 ;
	    RECT 6.2250 0.5300 6.6900 0.5800 ;
	    RECT 5.4450 0.3200 6.6900 0.5300 ;
	    RECT 7.0150 0.3700 7.3050 0.9200 ;
	    RECT 8.0250 0.7300 8.1950 2.3450 ;
	    RECT 7.8950 0.3200 8.1950 0.7300 ;
         LAYER met1 ;
	    RECT 2.8450 2.0000 3.1350 2.0550 ;
	    RECT 5.1450 2.0000 5.4350 2.0550 ;
	    RECT 2.8450 1.8250 5.4350 2.0000 ;
	    RECT 2.8450 1.7700 3.1350 1.8250 ;
	    RECT 5.1450 1.7700 5.4350 1.8250 ;
	    RECT 3.7650 1.1900 4.0550 1.2050 ;
	    RECT 5.1050 1.1900 5.4350 1.2050 ;
	    RECT 3.7650 1.1500 5.4350 1.1900 ;
	    RECT 6.5250 1.1500 6.8150 1.2050 ;
	    RECT 3.7650 0.9750 6.8150 1.1500 ;
	    RECT 3.7650 0.9600 5.4350 0.9750 ;
	    RECT 3.7650 0.9200 4.0550 0.9600 ;
	    RECT 5.1050 0.9200 5.4350 0.9600 ;
	    RECT 6.5250 0.9200 6.8150 0.9750 ;
	    RECT 4.2250 0.7250 4.5150 0.7800 ;
	    RECT 6.9850 0.7250 7.2750 0.7800 ;
	    RECT 4.2250 0.5500 7.2750 0.7250 ;
	    RECT 4.2250 0.4950 4.5150 0.5500 ;
	    RECT 6.9850 0.4950 7.2750 0.5500 ;
   END
END efs8hd_xnor3_1
MACRO efs8hd_xnor3_2
   CLASS CORE ;
   FOREIGN efs8hd_xnor3_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 8.7400 BY 3.4000 ;
   SITE unitehd ;
   PIN C
      PORT
         LAYER li1 ;
	    RECT 2.0750 1.3450 2.6400 1.6550 ;
      END
   END C
   PIN A
      PORT
         LAYER li1 ;
	    RECT 7.5050 1.3450 7.9150 1.6550 ;
      END
   END A
   PIN B
      PORT
         LAYER li1 ;
	    RECT 6.5850 1.7850 7.2650 2.0200 ;
	    RECT 6.5850 1.2450 6.8550 1.7850 ;
      END
   END B
   PIN X
      PORT
         LAYER li1 ;
	    RECT 0.5450 1.8000 0.8250 3.0800 ;
	    RECT 0.5450 1.1550 0.7900 1.8000 ;
	    RECT 0.5450 0.4400 0.8050 1.1550 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.1050 0.3750 0.9200 ;
	    RECT 0.9750 0.1050 1.2250 0.6550 ;
	    RECT 3.9350 0.1050 4.1050 1.0800 ;
	    RECT 7.9350 0.1050 8.1050 0.7050 ;
	    RECT 0.0850 0.0850 8.1050 0.1050 ;
	    RECT 0.0000 -0.0850 8.7400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 8.7400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 8.7400 3.4850 ;
	    RECT 0.0850 3.2950 8.1900 3.3150 ;
	    RECT 0.0850 1.8650 0.3750 3.2950 ;
	    RECT 0.9950 2.7700 1.3300 3.2950 ;
	    RECT 3.6850 2.7950 4.0150 3.2950 ;
	    RECT 7.8550 2.8450 8.1900 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 8.7400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 1.5100 2.7950 2.9800 3.0050 ;
	    RECT 4.3500 2.8450 7.4450 3.0550 ;
	    RECT 1.5100 2.5550 1.6800 2.7950 ;
	    RECT 4.3500 2.5800 4.5200 2.8450 ;
	    RECT 0.9950 2.3450 1.6800 2.5550 ;
	    RECT 2.0200 2.3700 4.5200 2.5800 ;
	    RECT 0.9950 1.6550 1.1650 2.3450 ;
	    RECT 1.3950 1.9200 2.9800 2.1300 ;
	    RECT 0.9600 1.2450 1.1650 1.6550 ;
	    RECT 0.9900 1.0800 1.1650 1.2450 ;
	    RECT 0.9900 0.8700 1.5650 1.0800 ;
	    RECT 1.3950 0.5300 1.5650 0.8700 ;
	    RECT 1.7350 0.7450 1.9050 1.9200 ;
	    RECT 2.8100 1.6550 2.9800 1.9200 ;
	    RECT 3.1500 1.9050 3.5350 2.1200 ;
	    RECT 3.2550 1.7200 3.5350 1.9050 ;
	    RECT 2.8100 1.2450 3.0850 1.6550 ;
	    RECT 2.2050 0.9950 2.5850 1.1300 ;
	    RECT 3.2550 0.9950 3.4250 1.7200 ;
	    RECT 3.7050 1.5050 3.8750 2.3700 ;
	    RECT 4.1050 1.8050 4.5250 2.1450 ;
	    RECT 2.2050 0.7800 3.4250 0.9950 ;
	    RECT 3.5950 1.2950 3.8750 1.5050 ;
	    RECT 3.5950 0.5700 3.7650 1.2950 ;
	    RECT 2.5300 0.5300 2.9650 0.5700 ;
	    RECT 1.3950 0.3200 2.9650 0.5300 ;
	    RECT 3.1350 0.3550 3.7650 0.5700 ;
	    RECT 4.2850 0.5200 4.5250 1.8050 ;
	    RECT 4.7050 0.7450 4.8750 2.6300 ;
	    RECT 5.0450 1.0750 5.2150 2.8450 ;
	    RECT 8.3600 2.6300 8.6550 3.0800 ;
	    RECT 5.3950 2.0200 5.8100 2.5550 ;
	    RECT 6.2450 2.4200 8.6550 2.6300 ;
	    RECT 5.3950 1.8050 6.0750 2.0200 ;
	    RECT 5.4100 1.2450 5.7350 1.5950 ;
	    RECT 5.0450 0.9000 5.3950 1.0750 ;
	    RECT 5.5650 0.9900 5.7350 1.2450 ;
	    RECT 5.0850 0.8550 5.3950 0.9000 ;
	    RECT 4.7050 0.5550 4.9150 0.7450 ;
	    RECT 5.0850 0.7250 5.4550 0.8550 ;
	    RECT 4.7050 0.3300 5.1150 0.5550 ;
	    RECT 5.2850 0.4000 5.4550 0.7250 ;
	    RECT 5.9050 0.5300 6.0750 1.8050 ;
	    RECT 6.2450 0.7450 6.4150 2.4200 ;
	    RECT 8.1700 2.3450 8.6550 2.4200 ;
	    RECT 7.4350 1.8700 8.2550 2.1300 ;
	    RECT 8.0850 1.6550 8.2550 1.8700 ;
	    RECT 7.0250 1.1800 7.3350 1.5950 ;
	    RECT 8.0850 1.2450 8.3150 1.6550 ;
	    RECT 7.0250 0.9150 7.2300 1.1800 ;
	    RECT 8.0850 1.1300 8.2550 1.2450 ;
	    RECT 7.5150 0.9400 8.2550 1.1300 ;
	    RECT 7.4750 0.9200 8.2550 0.9400 ;
	    RECT 6.6850 0.5300 7.1500 0.5800 ;
	    RECT 5.9050 0.3200 7.1500 0.5300 ;
	    RECT 7.4750 0.3700 7.7650 0.9200 ;
	    RECT 8.4850 0.7300 8.6550 2.3450 ;
	    RECT 8.3550 0.3200 8.6550 0.7300 ;
         LAYER met1 ;
	    RECT 3.3050 2.0000 3.5950 2.0550 ;
	    RECT 5.6050 2.0000 5.8950 2.0550 ;
	    RECT 3.3050 1.8250 5.8950 2.0000 ;
	    RECT 3.3050 1.7700 3.5950 1.8250 ;
	    RECT 5.6050 1.7700 5.8950 1.8250 ;
	    RECT 4.2250 1.1900 4.5150 1.2050 ;
	    RECT 5.5650 1.1900 5.8950 1.2050 ;
	    RECT 4.2250 1.1500 5.8950 1.1900 ;
	    RECT 6.9850 1.1500 7.2750 1.2050 ;
	    RECT 4.2250 0.9750 7.2750 1.1500 ;
	    RECT 4.2250 0.9600 5.8950 0.9750 ;
	    RECT 4.2250 0.9200 4.5150 0.9600 ;
	    RECT 5.5650 0.9200 5.8950 0.9600 ;
	    RECT 6.9850 0.9200 7.2750 0.9750 ;
	    RECT 4.6850 0.7250 4.9750 0.7800 ;
	    RECT 7.4450 0.7250 7.7350 0.7800 ;
	    RECT 4.6850 0.5500 7.7350 0.7250 ;
	    RECT 4.6850 0.4950 4.9750 0.5500 ;
	    RECT 7.4450 0.4950 7.7350 0.5500 ;
   END
END efs8hd_xnor3_2
MACRO efs8hd_xnor3_4
   CLASS CORE ;
   FOREIGN efs8hd_xnor3_4 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 9.6600 BY 3.4000 ;
   SITE unitehd ;
   PIN C
      PORT
         LAYER li1 ;
	    RECT 2.9050 1.3450 3.5600 1.6550 ;
      END
   END C
   PIN A
      PORT
         LAYER li1 ;
	    RECT 8.4250 1.3450 8.8350 1.6550 ;
      END
   END A
   PIN B
      PORT
         LAYER li1 ;
	    RECT 7.5050 1.7850 8.1850 2.0200 ;
	    RECT 7.5050 1.2450 7.7750 1.7850 ;
      END
   END B
   PIN X
      PORT
         LAYER li1 ;
	    RECT 0.6250 1.6550 0.9550 3.0300 ;
	    RECT 1.4650 1.8000 1.7450 3.0800 ;
	    RECT 1.4650 1.6550 1.7100 1.8000 ;
	    RECT 0.6250 1.2450 1.7100 1.6550 ;
	    RECT 0.6250 0.4700 0.8750 1.2450 ;
	    RECT 1.4650 1.1550 1.7100 1.2450 ;
	    RECT 1.4650 0.4400 1.7150 1.1550 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.2050 0.1050 0.4550 0.9200 ;
	    RECT 1.0450 0.1050 1.2950 0.9200 ;
	    RECT 1.8850 0.1050 2.0550 0.6550 ;
	    RECT 4.8550 0.1050 5.0250 1.0800 ;
	    RECT 8.8550 0.1050 9.0250 0.7050 ;
	    RECT 0.2050 0.0850 9.0250 0.1050 ;
	    RECT 0.0000 -0.0850 9.6600 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 9.6600 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 9.6600 3.4850 ;
	    RECT 0.2050 3.2950 9.1100 3.3150 ;
	    RECT 0.2050 1.8650 0.4550 3.2950 ;
	    RECT 1.1250 1.8700 1.2950 3.2950 ;
	    RECT 1.9150 2.7700 2.2500 3.2950 ;
	    RECT 4.6050 2.7950 4.9350 3.2950 ;
	    RECT 8.7750 2.8450 9.1100 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 9.6600 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 2.4300 2.7950 3.9000 3.0050 ;
	    RECT 5.2700 2.8450 8.3650 3.0550 ;
	    RECT 2.4300 2.5550 2.6000 2.7950 ;
	    RECT 5.2700 2.5800 5.4400 2.8450 ;
	    RECT 1.9150 2.3450 2.6000 2.5550 ;
	    RECT 2.9400 2.3700 5.4400 2.5800 ;
	    RECT 1.9150 1.6550 2.0850 2.3450 ;
	    RECT 2.3150 1.9200 3.9000 2.1300 ;
	    RECT 1.8800 1.2450 2.0850 1.6550 ;
	    RECT 1.9100 1.0800 2.0850 1.2450 ;
	    RECT 1.9100 0.8700 2.3950 1.0800 ;
	    RECT 2.2250 0.5300 2.3950 0.8700 ;
	    RECT 2.5650 0.7450 2.7350 1.9200 ;
	    RECT 3.7300 1.6550 3.9000 1.9200 ;
	    RECT 4.0700 1.9050 4.4550 2.1200 ;
	    RECT 4.1750 1.7200 4.4550 1.9050 ;
	    RECT 3.7300 1.2450 4.0050 1.6550 ;
	    RECT 3.1250 0.9950 3.5050 1.1300 ;
	    RECT 4.1750 0.9950 4.3450 1.7200 ;
	    RECT 4.6250 1.5050 4.7950 2.3700 ;
	    RECT 5.0250 1.8050 5.4450 2.1450 ;
	    RECT 3.1250 0.7800 4.3450 0.9950 ;
	    RECT 4.5150 1.2950 4.7950 1.5050 ;
	    RECT 4.5150 0.5700 4.6850 1.2950 ;
	    RECT 3.4500 0.5300 3.8850 0.5700 ;
	    RECT 2.2250 0.3200 3.8850 0.5300 ;
	    RECT 4.0550 0.3550 4.6850 0.5700 ;
	    RECT 5.2050 0.5200 5.4450 1.8050 ;
	    RECT 5.6250 0.7450 5.7950 2.6300 ;
	    RECT 5.9650 1.0750 6.1350 2.8450 ;
	    RECT 9.2800 2.6300 9.5750 3.0800 ;
	    RECT 6.3150 2.0200 6.7300 2.5550 ;
	    RECT 7.1650 2.4200 9.5750 2.6300 ;
	    RECT 6.3150 1.8050 6.9950 2.0200 ;
	    RECT 6.3300 1.2450 6.6550 1.5950 ;
	    RECT 5.9650 0.9000 6.3150 1.0750 ;
	    RECT 6.4850 0.9900 6.6550 1.2450 ;
	    RECT 6.0050 0.8550 6.3150 0.9000 ;
	    RECT 5.6250 0.5550 5.8350 0.7450 ;
	    RECT 6.0050 0.7250 6.3750 0.8550 ;
	    RECT 5.6250 0.3300 6.0350 0.5550 ;
	    RECT 6.2050 0.4000 6.3750 0.7250 ;
	    RECT 6.8250 0.5300 6.9950 1.8050 ;
	    RECT 7.1650 0.7450 7.3350 2.4200 ;
	    RECT 9.0900 2.3450 9.5750 2.4200 ;
	    RECT 8.3550 1.8700 9.1750 2.1300 ;
	    RECT 9.0050 1.6550 9.1750 1.8700 ;
	    RECT 7.9450 1.1800 8.2550 1.5950 ;
	    RECT 9.0050 1.2450 9.2350 1.6550 ;
	    RECT 7.9450 0.9150 8.1500 1.1800 ;
	    RECT 9.0050 1.1300 9.1750 1.2450 ;
	    RECT 8.4350 0.9400 9.1750 1.1300 ;
	    RECT 8.3950 0.9200 9.1750 0.9400 ;
	    RECT 7.6050 0.5300 8.0700 0.5800 ;
	    RECT 6.8250 0.3200 8.0700 0.5300 ;
	    RECT 8.3950 0.3700 8.6850 0.9200 ;
	    RECT 9.4050 0.7300 9.5750 2.3450 ;
	    RECT 9.2750 0.3200 9.5750 0.7300 ;
         LAYER met1 ;
	    RECT 4.2250 2.0000 4.5150 2.0550 ;
	    RECT 6.5250 2.0000 6.8150 2.0550 ;
	    RECT 4.2250 1.8250 6.8150 2.0000 ;
	    RECT 4.2250 1.7700 4.5150 1.8250 ;
	    RECT 6.5250 1.7700 6.8150 1.8250 ;
	    RECT 5.1450 1.1900 5.4350 1.2050 ;
	    RECT 6.4850 1.1900 6.8150 1.2050 ;
	    RECT 5.1450 1.1500 6.8150 1.1900 ;
	    RECT 7.9050 1.1500 8.1950 1.2050 ;
	    RECT 5.1450 0.9750 8.1950 1.1500 ;
	    RECT 5.1450 0.9600 6.8150 0.9750 ;
	    RECT 5.1450 0.9200 5.4350 0.9600 ;
	    RECT 6.4850 0.9200 6.8150 0.9600 ;
	    RECT 7.9050 0.9200 8.1950 0.9750 ;
	    RECT 5.6050 0.7250 5.8950 0.7800 ;
	    RECT 8.3650 0.7250 8.6550 0.7800 ;
	    RECT 5.6050 0.5500 8.6550 0.7250 ;
	    RECT 5.6050 0.4950 5.8950 0.5500 ;
	    RECT 8.3650 0.4950 8.6550 0.5500 ;
   END
END efs8hd_xnor3_4
MACRO efs8hd_xor2_2
   CLASS CORE ;
   FOREIGN efs8hd_xor2_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 5.9800 BY 3.4000 ;
   SITE unitehd ;
   PIN B
      PORT
         LAYER li1 ;
	    RECT 1.0450 1.3450 1.5400 1.5950 ;
	    RECT 3.3650 1.3450 4.0900 1.6150 ;
         LAYER met1 ;
	    RECT 1.0050 1.5750 1.2950 1.6300 ;
	    RECT 3.7650 1.5750 4.0550 1.6300 ;
	    RECT 1.0050 1.4000 4.0550 1.5750 ;
	    RECT 1.0050 1.3450 1.2950 1.4000 ;
	    RECT 3.7650 1.3450 4.0550 1.4000 ;
      END
   END B
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.7050 1.8050 1.8800 2.0200 ;
	    RECT 0.7050 1.5950 0.8750 1.8050 ;
	    RECT 0.5450 1.3450 0.8750 1.5950 ;
	    RECT 1.7100 1.6300 1.8800 1.8050 ;
	    RECT 1.7100 1.3000 3.1950 1.6300 ;
      END
   END A
   PIN X
      PORT
         LAYER li1 ;
	    RECT 5.0250 2.0300 5.2750 2.6550 ;
	    RECT 5.0250 1.7700 5.8950 2.0300 ;
	    RECT 5.4850 1.1300 5.8950 1.7700 ;
	    RECT 3.6250 0.9050 5.8950 1.1300 ;
	    RECT 3.6250 0.8050 3.9550 0.9050 ;
	    RECT 4.9850 0.8050 5.3150 0.9050 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1900 0.1050 0.3600 0.6950 ;
	    RECT 1.0300 0.1050 1.2000 0.6950 ;
	    RECT 1.8700 0.1050 2.0400 0.6950 ;
	    RECT 2.8100 0.1050 2.9800 0.6950 ;
	    RECT 4.6450 0.1050 4.8150 0.6950 ;
	    RECT 5.4850 0.1050 5.6550 0.6950 ;
	    RECT 0.1900 0.0850 5.6550 0.1050 ;
	    RECT 0.0000 -0.0850 5.9800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 5.9800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 5.9800 3.4850 ;
	    RECT 0.5700 3.2950 3.9150 3.3150 ;
	    RECT 0.5700 2.6700 0.8200 3.2950 ;
	    RECT 2.7700 2.6700 3.0200 3.2950 ;
	    RECT 3.6100 2.6700 3.9150 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 5.9800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.1200 2.6700 0.4000 3.0800 ;
	    RECT 0.9900 2.8700 2.0800 3.0800 ;
	    RECT 0.9900 2.6700 1.2400 2.8700 ;
	    RECT 1.8300 2.6700 2.0800 2.8700 ;
	    RECT 0.1450 2.6550 0.3150 2.6700 ;
	    RECT 1.0650 2.6550 1.2350 2.6700 ;
	    RECT 2.2850 2.6550 2.6000 3.0800 ;
	    RECT 1.4100 2.4450 1.6600 2.6550 ;
	    RECT 2.3900 2.4450 2.6000 2.6550 ;
	    RECT 3.1900 2.4450 3.4400 3.0800 ;
	    RECT 4.0850 2.8700 5.6950 3.0800 ;
	    RECT 4.0850 2.4450 4.8550 2.8700 ;
	    RECT 0.1200 2.2300 2.2200 2.4450 ;
	    RECT 2.3900 2.2300 4.8550 2.4450 ;
	    RECT 5.4450 2.2450 5.6950 2.8700 ;
	    RECT 0.1200 1.1300 0.2900 2.2300 ;
	    RECT 2.0500 2.0200 2.2200 2.2300 ;
	    RECT 2.0500 1.8050 4.7850 2.0200 ;
	    RECT 4.6150 1.5550 4.7850 1.8050 ;
	    RECT 4.6150 1.3450 5.2750 1.5550 ;
	    RECT 0.1200 0.9050 1.7000 1.1300 ;
	    RECT 0.5300 0.3200 0.8600 0.9050 ;
	    RECT 1.3700 0.3200 1.7000 0.9050 ;
	    RECT 2.3100 0.9050 3.4000 1.1300 ;
	    RECT 2.3100 0.3200 2.6400 0.9050 ;
	    RECT 3.1500 0.5950 3.4000 0.9050 ;
	    RECT 3.1500 0.3200 4.3800 0.5950 ;
         LAYER met1 ;
	    RECT 0.0850 2.8500 0.3750 2.9050 ;
	    RECT 1.0050 2.8500 1.2950 2.9050 ;
	    RECT 0.0850 2.6750 1.2950 2.8500 ;
	    RECT 0.0850 2.6200 0.3750 2.6750 ;
	    RECT 1.0050 2.6200 1.2950 2.6750 ;
   END
END efs8hd_xor2_2
MACRO efs8hd_xor2_4
   CLASS CORE ;
   FOREIGN efs8hd_xor2_4 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 10.1200 BY 3.4000 ;
   SITE unitehd ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 2.6300 1.7850 6.1650 2.0200 ;
	    RECT 2.6300 1.5950 2.8000 1.7850 ;
	    RECT 0.4250 1.3450 2.8000 1.5950 ;
	    RECT 5.9950 1.5950 6.1650 1.7850 ;
	    RECT 5.9950 1.3450 7.3700 1.5950 ;
      END
   END A
   PIN B
      PORT
         LAYER li1 ;
	    RECT 2.9700 1.3800 5.7400 1.6150 ;
	    RECT 2.9700 1.3450 5.0000 1.3800 ;
      END
   END B
   PIN X
      PORT
         LAYER li1 ;
	    RECT 7.8800 2.0800 8.1700 2.6550 ;
	    RECT 8.7600 2.0800 9.0100 2.6550 ;
	    RECT 7.8800 2.0300 9.0100 2.0800 ;
	    RECT 9.6000 2.0300 10.0350 3.0800 ;
	    RECT 7.8800 1.8050 10.0350 2.0300 ;
	    RECT 5.1500 1.1300 5.5800 1.1700 ;
	    RECT 4.1650 0.8050 5.5800 1.1300 ;
	    RECT 7.8500 1.1300 8.3050 1.1700 ;
	    RECT 9.7350 1.1300 10.0350 1.8050 ;
	    RECT 7.8500 0.9200 10.0350 1.1300 ;
	    RECT 7.8500 0.9050 8.6300 0.9200 ;
	    RECT 8.3000 0.3200 8.6300 0.9050 ;
	    RECT 9.1400 0.3200 9.4700 0.9200 ;
         LAYER met1 ;
	    RECT 5.1450 1.1500 5.4350 1.2050 ;
	    RECT 7.9050 1.1500 8.1950 1.2050 ;
	    RECT 5.1450 0.9750 8.1950 1.1500 ;
	    RECT 5.1450 0.9200 5.4350 0.9750 ;
	    RECT 7.9050 0.9200 8.1950 0.9750 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.0850 0.1050 0.3600 0.7050 ;
	    RECT 1.0300 0.1050 1.2000 0.6950 ;
	    RECT 1.8700 0.1050 2.0400 0.6950 ;
	    RECT 2.7100 0.1050 2.8800 0.6950 ;
	    RECT 3.5500 0.1050 3.8200 1.1200 ;
	    RECT 6.1700 0.1050 6.3400 0.6950 ;
	    RECT 7.0100 0.1050 7.1800 0.6950 ;
	    RECT 7.9600 0.1050 8.1300 0.6950 ;
	    RECT 8.8000 0.1050 8.9700 0.6950 ;
	    RECT 9.6400 0.1050 9.8100 0.6950 ;
	    RECT 0.0850 0.0850 9.8100 0.1050 ;
	    RECT 0.0000 -0.0850 10.1200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 10.1200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 10.1200 3.4850 ;
	    RECT 0.5700 3.2950 7.2200 3.3150 ;
	    RECT 0.5700 2.7200 0.8200 3.2950 ;
	    RECT 1.4100 2.7200 1.6600 3.2950 ;
	    RECT 4.4500 2.7200 4.7000 3.2950 ;
	    RECT 5.2900 2.7200 5.5400 3.2950 ;
	    RECT 6.1300 2.7200 6.3800 3.2950 ;
	    RECT 6.9700 2.7200 7.2200 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 10.1200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 0.0850 2.5050 0.4000 3.0800 ;
	    RECT 0.9900 2.5050 1.2400 3.0800 ;
	    RECT 1.8300 2.8700 3.7600 3.0800 ;
	    RECT 1.8300 2.5050 2.0800 2.8700 ;
	    RECT 2.6700 2.6550 2.9200 2.8700 ;
	    RECT 0.0850 2.2300 2.0800 2.5050 ;
	    RECT 2.2500 2.4450 2.5000 2.6550 ;
	    RECT 3.0900 2.4450 3.3400 2.6550 ;
	    RECT 2.2500 2.2300 3.3400 2.4450 ;
	    RECT 3.5100 2.2450 3.7600 2.8700 ;
	    RECT 4.0300 2.5050 4.2800 3.0800 ;
	    RECT 4.8700 2.5050 5.1200 3.0800 ;
	    RECT 5.7100 2.5050 5.9600 3.0800 ;
	    RECT 6.5500 2.5050 6.8000 3.0800 ;
	    RECT 7.3900 2.8700 9.4300 3.0800 ;
	    RECT 7.3900 2.5050 7.6400 2.8700 ;
	    RECT 4.0300 2.2300 7.6400 2.5050 ;
	    RECT 8.3400 2.2950 8.5900 2.8700 ;
	    RECT 9.1800 2.2450 9.4300 2.8700 ;
	    RECT 2.2500 2.0200 2.4200 2.2300 ;
	    RECT 0.0850 1.8050 2.4200 2.0200 ;
	    RECT 6.5500 1.8200 6.8000 2.2300 ;
	    RECT 7.2600 1.8050 7.7100 2.0200 ;
	    RECT 0.0850 1.1300 0.2550 1.8050 ;
	    RECT 7.5400 1.5950 7.7100 1.8050 ;
	    RECT 7.5400 1.3800 9.5650 1.5950 ;
	    RECT 8.5400 1.3450 9.5650 1.3800 ;
	    RECT 0.0850 0.9200 3.3800 1.1300 ;
	    RECT 0.5300 0.9050 3.3800 0.9200 ;
	    RECT 0.5300 0.3200 0.8600 0.9050 ;
	    RECT 1.3700 0.3200 1.7000 0.9050 ;
	    RECT 2.2100 0.3200 2.5400 0.9050 ;
	    RECT 3.0500 0.3200 3.3800 0.9050 ;
	    RECT 5.7500 0.9050 7.6800 1.1300 ;
	    RECT 5.7500 0.5950 6.0000 0.9050 ;
	    RECT 3.9900 0.3200 6.0000 0.5950 ;
	    RECT 6.5100 0.3200 6.8400 0.9050 ;
	    RECT 7.3500 0.3200 7.6800 0.9050 ;
         LAYER met1 ;
	    RECT 1.9250 2.0000 2.2150 2.0550 ;
	    RECT 7.4450 2.0000 7.7350 2.0550 ;
	    RECT 1.9250 1.8250 7.7350 2.0000 ;
	    RECT 1.9250 1.7700 2.2150 1.8250 ;
	    RECT 7.4450 1.7700 7.7350 1.8250 ;
   END
END efs8hd_xor2_4
MACRO efs8hd_xor3_1
   CLASS CORE ;
   FOREIGN efs8hd_xor3_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 8.7400 BY 3.4000 ;
   SITE unitehd ;
   PIN C
      PORT
         LAYER li1 ;
	    RECT 1.8600 1.1050 2.6150 1.6550 ;
      END
   END C
   PIN A
      PORT
         LAYER li1 ;
	    RECT 7.5050 1.3450 7.9150 1.6550 ;
      END
   END A
   PIN B
      PORT
         LAYER li1 ;
	    RECT 6.5850 1.7850 7.2650 2.0200 ;
	    RECT 6.5850 1.2450 6.8550 1.7850 ;
      END
   END B
   PIN X
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.8000 0.6100 3.0800 ;
	    RECT 0.0850 1.1550 0.4000 1.8000 ;
	    RECT 0.0850 0.4400 0.5900 1.1550 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.7600 0.1050 1.0100 0.6550 ;
	    RECT 3.9300 0.1050 4.1000 1.0800 ;
	    RECT 7.9350 0.1050 8.1050 0.7050 ;
	    RECT 0.7600 0.0850 8.1050 0.1050 ;
	    RECT 0.0000 -0.0850 8.7400 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 8.7400 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 8.7400 3.4850 ;
	    RECT 0.7800 3.2950 8.1900 3.3150 ;
	    RECT 0.7800 2.7700 1.1150 3.2950 ;
	    RECT 3.8050 2.7550 4.0150 3.2950 ;
	    RECT 7.8550 2.8450 8.1900 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 8.7400 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 1.3000 2.7950 2.8950 3.0050 ;
	    RECT 3.1100 2.7950 3.6350 3.0050 ;
	    RECT 1.3000 2.5550 1.4700 2.7950 ;
	    RECT 3.4650 2.5800 3.6350 2.7950 ;
	    RECT 4.3500 2.8450 7.4450 3.0550 ;
	    RECT 4.3500 2.5800 4.5200 2.8450 ;
	    RECT 0.7800 2.3450 1.4700 2.5550 ;
	    RECT 1.8700 2.3700 3.2950 2.5800 ;
	    RECT 3.4650 2.3700 4.5200 2.5800 ;
	    RECT 0.7800 1.6550 0.9500 2.3450 ;
	    RECT 1.1850 1.9200 2.9550 2.1300 ;
	    RECT 0.7500 1.2450 0.9500 1.6550 ;
	    RECT 0.7800 1.0800 0.9500 1.2450 ;
	    RECT 0.7800 0.8700 1.3500 1.0800 ;
	    RECT 1.1800 0.5300 1.3500 0.8700 ;
	    RECT 1.5200 0.7450 1.6900 1.9200 ;
	    RECT 2.7850 1.2450 2.9550 1.9200 ;
	    RECT 3.1250 2.1200 3.2950 2.3700 ;
	    RECT 3.1250 1.9050 3.5350 2.1200 ;
	    RECT 3.2500 1.7200 3.5350 1.9050 ;
	    RECT 1.9700 0.7650 3.0800 0.9350 ;
	    RECT 2.3900 0.5300 2.7400 0.5700 ;
	    RECT 1.1800 0.3200 2.7400 0.5300 ;
	    RECT 2.9100 0.5300 3.0800 0.7650 ;
	    RECT 3.2500 0.7450 3.4200 1.7200 ;
	    RECT 3.7050 1.5050 3.8750 2.3700 ;
	    RECT 4.1050 1.8050 4.5200 2.1450 ;
	    RECT 3.5900 1.2950 3.8750 1.5050 ;
	    RECT 3.5900 0.5300 3.7600 1.2950 ;
	    RECT 2.9100 0.3200 3.7600 0.5300 ;
	    RECT 4.2800 0.5200 4.5200 1.8050 ;
	    RECT 4.6950 0.7450 4.9050 2.6300 ;
	    RECT 5.0750 1.0750 5.2450 2.8450 ;
	    RECT 8.3600 2.6300 8.6550 3.0800 ;
	    RECT 5.4150 2.0200 5.8100 2.5550 ;
	    RECT 6.2450 2.4200 8.6550 2.6300 ;
	    RECT 5.4150 1.8050 6.0750 2.0200 ;
	    RECT 5.4150 1.2450 5.7350 1.5950 ;
	    RECT 5.0750 0.9000 5.3950 1.0750 ;
	    RECT 5.5650 0.9900 5.7350 1.2450 ;
	    RECT 5.0850 0.8600 5.3950 0.9000 ;
	    RECT 4.6950 0.5650 4.9150 0.7450 ;
	    RECT 5.0850 0.7350 5.4500 0.8600 ;
	    RECT 4.6950 0.3300 5.1100 0.5650 ;
	    RECT 5.2800 0.4000 5.4500 0.7350 ;
	    RECT 5.9050 0.5300 6.0750 1.8050 ;
	    RECT 6.2450 0.7450 6.4150 2.4200 ;
	    RECT 8.1700 2.3450 8.6550 2.4200 ;
	    RECT 7.4350 1.8700 8.2550 2.1300 ;
	    RECT 8.0850 1.6550 8.2550 1.8700 ;
	    RECT 7.0250 1.1800 7.3350 1.5950 ;
	    RECT 8.0850 1.2450 8.3150 1.6550 ;
	    RECT 7.0250 0.9150 7.2300 1.1800 ;
	    RECT 8.0850 1.1300 8.2550 1.2450 ;
	    RECT 7.5150 0.9400 8.2550 1.1300 ;
	    RECT 7.4750 0.9200 8.2550 0.9400 ;
	    RECT 6.6850 0.5300 7.1500 0.5800 ;
	    RECT 5.9050 0.3200 7.1500 0.5300 ;
	    RECT 7.4750 0.3700 7.7650 0.9200 ;
	    RECT 8.4850 0.7300 8.6550 2.3450 ;
	    RECT 8.3550 0.3200 8.6550 0.7300 ;
         LAYER met1 ;
	    RECT 3.3050 2.0000 3.5950 2.0550 ;
	    RECT 5.6050 2.0000 5.8950 2.0550 ;
	    RECT 3.3050 1.8250 5.8950 2.0000 ;
	    RECT 3.3050 1.7700 3.5950 1.8250 ;
	    RECT 5.6050 1.7700 5.8950 1.8250 ;
	    RECT 4.2250 1.1900 4.5150 1.2050 ;
	    RECT 5.5650 1.1900 5.8950 1.2050 ;
	    RECT 4.2250 1.1500 5.8950 1.1900 ;
	    RECT 6.9850 1.1500 7.2750 1.2050 ;
	    RECT 4.2250 0.9750 7.2750 1.1500 ;
	    RECT 4.2250 0.9600 5.8950 0.9750 ;
	    RECT 4.2250 0.9200 4.5150 0.9600 ;
	    RECT 5.5650 0.9200 5.8950 0.9600 ;
	    RECT 6.9850 0.9200 7.2750 0.9750 ;
	    RECT 4.6850 0.7250 4.9750 0.7800 ;
	    RECT 7.4450 0.7250 7.7350 0.7800 ;
	    RECT 4.6850 0.5500 7.7350 0.7250 ;
	    RECT 4.6850 0.4950 4.9750 0.5500 ;
	    RECT 7.4450 0.4950 7.7350 0.5500 ;
   END
END efs8hd_xor3_1
MACRO efs8hd_xor3_2
   CLASS CORE ;
   FOREIGN efs8hd_xor3_2 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 9.2000 BY 3.4000 ;
   SITE unitehd ;
   PIN C
      PORT
         LAYER li1 ;
	    RECT 2.3200 1.1050 3.0750 1.6550 ;
      END
   END C
   PIN A
      PORT
         LAYER li1 ;
	    RECT 7.9650 1.3450 8.3750 1.6550 ;
      END
   END A
   PIN B
      PORT
         LAYER li1 ;
	    RECT 7.0450 1.7850 7.7250 2.0200 ;
	    RECT 7.0450 1.2450 7.3150 1.7850 ;
      END
   END B
   PIN X
      PORT
         LAYER li1 ;
	    RECT 0.8200 2.5550 1.0700 3.0800 ;
	    RECT 0.5450 1.8000 1.0700 2.5550 ;
	    RECT 0.5450 1.1550 0.8600 1.8000 ;
	    RECT 0.5450 0.8250 1.0500 1.1550 ;
	    RECT 0.8000 0.4400 1.0500 0.8250 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.3000 0.1050 0.6300 0.5800 ;
	    RECT 1.2200 0.1050 1.4700 0.6550 ;
	    RECT 4.3900 0.1050 4.5600 1.0800 ;
	    RECT 8.3950 0.1050 8.5650 0.7050 ;
	    RECT 0.3000 0.0850 8.5650 0.1050 ;
	    RECT 0.0000 -0.0850 9.2000 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 9.2000 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 9.2000 3.4850 ;
	    RECT 0.3000 3.2950 8.6500 3.3150 ;
	    RECT 0.3000 2.7700 0.6500 3.2950 ;
	    RECT 1.2400 2.7700 1.5750 3.2950 ;
	    RECT 4.2650 2.7550 4.4750 3.2950 ;
	    RECT 8.3150 2.8450 8.6500 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 9.2000 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 1.7600 2.7950 3.3550 3.0050 ;
	    RECT 3.5700 2.7950 4.0950 3.0050 ;
	    RECT 1.7600 2.5550 1.9300 2.7950 ;
	    RECT 3.9250 2.5800 4.0950 2.7950 ;
	    RECT 4.8100 2.8450 7.9050 3.0550 ;
	    RECT 4.8100 2.5800 4.9800 2.8450 ;
	    RECT 1.2400 2.3450 1.9300 2.5550 ;
	    RECT 2.3300 2.3700 3.7550 2.5800 ;
	    RECT 3.9250 2.3700 4.9800 2.5800 ;
	    RECT 1.2400 1.6550 1.4100 2.3450 ;
	    RECT 1.6450 1.9200 3.4150 2.1300 ;
	    RECT 1.2100 1.2450 1.4100 1.6550 ;
	    RECT 1.2400 1.0800 1.4100 1.2450 ;
	    RECT 1.2400 0.8700 1.8100 1.0800 ;
	    RECT 1.6400 0.5300 1.8100 0.8700 ;
	    RECT 1.9800 0.7450 2.1500 1.9200 ;
	    RECT 3.2450 1.2450 3.4150 1.9200 ;
	    RECT 3.5850 2.1200 3.7550 2.3700 ;
	    RECT 3.5850 1.9050 3.9950 2.1200 ;
	    RECT 3.7100 1.7200 3.9950 1.9050 ;
	    RECT 2.4300 0.7650 3.5400 0.9350 ;
	    RECT 2.8500 0.5300 3.2000 0.5700 ;
	    RECT 1.6400 0.3200 3.2000 0.5300 ;
	    RECT 3.3700 0.5300 3.5400 0.7650 ;
	    RECT 3.7100 0.7450 3.8800 1.7200 ;
	    RECT 4.1650 1.5050 4.3350 2.3700 ;
	    RECT 4.5650 1.8050 4.9800 2.1450 ;
	    RECT 4.0500 1.2950 4.3350 1.5050 ;
	    RECT 4.0500 0.5300 4.2200 1.2950 ;
	    RECT 3.3700 0.3200 4.2200 0.5300 ;
	    RECT 4.7400 0.5200 4.9800 1.8050 ;
	    RECT 5.1550 0.7450 5.3650 2.6300 ;
	    RECT 5.5350 1.0750 5.7050 2.8450 ;
	    RECT 8.8200 2.6300 9.1150 3.0800 ;
	    RECT 5.8750 2.0200 6.2700 2.5550 ;
	    RECT 6.7050 2.4200 9.1150 2.6300 ;
	    RECT 5.8750 1.8050 6.5350 2.0200 ;
	    RECT 5.8750 1.2450 6.1950 1.5950 ;
	    RECT 5.5350 0.9000 5.8550 1.0750 ;
	    RECT 6.0250 0.9900 6.1950 1.2450 ;
	    RECT 5.5450 0.8600 5.8550 0.9000 ;
	    RECT 5.1550 0.5650 5.3750 0.7450 ;
	    RECT 5.5450 0.7350 5.9100 0.8600 ;
	    RECT 5.1550 0.3300 5.5700 0.5650 ;
	    RECT 5.7400 0.4000 5.9100 0.7350 ;
	    RECT 6.3650 0.5300 6.5350 1.8050 ;
	    RECT 6.7050 0.7450 6.8750 2.4200 ;
	    RECT 8.6300 2.3450 9.1150 2.4200 ;
	    RECT 7.8950 1.8700 8.7150 2.1300 ;
	    RECT 8.5450 1.6550 8.7150 1.8700 ;
	    RECT 7.4850 1.1800 7.7950 1.5950 ;
	    RECT 8.5450 1.2450 8.7750 1.6550 ;
	    RECT 7.4850 0.9150 7.6900 1.1800 ;
	    RECT 8.5450 1.1300 8.7150 1.2450 ;
	    RECT 7.9750 0.9400 8.7150 1.1300 ;
	    RECT 7.9350 0.9200 8.7150 0.9400 ;
	    RECT 7.1450 0.5300 7.6100 0.5800 ;
	    RECT 6.3650 0.3200 7.6100 0.5300 ;
	    RECT 7.9350 0.3700 8.2250 0.9200 ;
	    RECT 8.9450 0.7300 9.1150 2.3450 ;
	    RECT 8.8150 0.3200 9.1150 0.7300 ;
         LAYER met1 ;
	    RECT 3.7650 2.0000 4.0550 2.0550 ;
	    RECT 6.0650 2.0000 6.3550 2.0550 ;
	    RECT 3.7650 1.8250 6.3550 2.0000 ;
	    RECT 3.7650 1.7700 4.0550 1.8250 ;
	    RECT 6.0650 1.7700 6.3550 1.8250 ;
	    RECT 4.6850 1.2000 4.9750 1.2050 ;
	    RECT 6.0250 1.2000 6.3550 1.2050 ;
	    RECT 4.6850 1.1500 6.3550 1.2000 ;
	    RECT 7.4450 1.1500 7.7350 1.2050 ;
	    RECT 4.6850 0.9750 7.7350 1.1500 ;
	    RECT 4.6850 0.9700 6.3550 0.9750 ;
	    RECT 4.6850 0.9200 4.9750 0.9700 ;
	    RECT 6.0250 0.9200 6.3550 0.9700 ;
	    RECT 7.4450 0.9200 7.7350 0.9750 ;
	    RECT 5.1450 0.7250 5.4350 0.7800 ;
	    RECT 7.9050 0.7250 8.1950 0.7800 ;
	    RECT 5.1450 0.5500 8.1950 0.7250 ;
	    RECT 5.1450 0.4950 5.4350 0.5500 ;
	    RECT 7.9050 0.4950 8.1950 0.5500 ;
   END
END efs8hd_xor3_2
MACRO efs8hd_xor3_4
   CLASS CORE ;
   FOREIGN efs8hd_xor3_4 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 10.1200 BY 3.4000 ;
   SITE unitehd ;
   PIN C
      PORT
         LAYER li1 ;
	    RECT 2.8800 1.1050 3.5350 1.6550 ;
      END
   END C
   PIN A
      PORT
         LAYER li1 ;
	    RECT 8.4250 1.3450 9.0550 1.6550 ;
      END
   END A
   PIN B
      PORT
         LAYER li1 ;
	    RECT 7.5050 1.7850 8.2850 2.0200 ;
	    RECT 7.5050 1.2450 7.8750 1.7850 ;
      END
   END B
   PIN X
      PORT
         LAYER li1 ;
	    RECT 0.6950 2.5550 0.8650 3.0800 ;
	    RECT 1.5350 2.5550 1.7050 3.0800 ;
	    RECT 0.6950 1.8200 1.7050 2.5550 ;
	    RECT 0.6950 1.7850 1.4200 1.8200 ;
	    RECT 1.1050 1.1550 1.4200 1.7850 ;
	    RECT 0.5950 1.0400 1.5350 1.1550 ;
	    RECT 0.5950 0.8250 1.6050 1.0400 ;
	    RECT 0.5950 0.4400 0.7650 0.8250 ;
	    RECT 1.4350 0.4400 1.6050 0.8250 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.1750 0.1050 0.3450 0.6800 ;
	    RECT 0.9350 0.1050 1.2650 0.5800 ;
	    RECT 1.8550 0.1050 2.0250 0.6550 ;
	    RECT 0.1750 0.0950 2.0250 0.1050 ;
	    RECT 4.8800 0.1050 5.1200 1.1050 ;
	    RECT 8.9950 0.1050 9.1650 0.7050 ;
	    RECT 4.8800 0.0950 9.1650 0.1050 ;
	    RECT 0.1750 0.0850 9.1650 0.0950 ;
	    RECT 0.0000 -0.0850 10.1200 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 10.1200 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 10.1200 3.4850 ;
	    RECT 0.2750 3.2950 9.2450 3.3150 ;
	    RECT 0.2750 2.6700 0.4450 3.2950 ;
	    RECT 1.0350 2.7700 1.3650 3.2950 ;
	    RECT 1.8750 2.7700 2.2050 3.2950 ;
	    RECT 4.7250 2.7550 5.0350 3.2950 ;
	    RECT 8.9150 2.8450 9.2450 3.2950 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 10.1200 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 2.3750 2.7950 3.9150 3.0050 ;
	    RECT 4.1300 2.7950 4.5550 3.0050 ;
	    RECT 2.3750 2.5550 2.5450 2.7950 ;
	    RECT 4.3850 2.5800 4.5550 2.7950 ;
	    RECT 5.3700 2.8450 8.4650 3.0550 ;
	    RECT 5.3700 2.5800 5.5400 2.8450 ;
	    RECT 1.8750 2.3450 2.5450 2.5550 ;
	    RECT 2.8900 2.3700 4.2150 2.5800 ;
	    RECT 4.3850 2.3700 5.5400 2.5800 ;
	    RECT 1.8750 1.6550 2.0450 2.3450 ;
	    RECT 2.3700 1.9200 3.8750 2.1300 ;
	    RECT 1.8200 1.2050 2.0450 1.6550 ;
	    RECT 1.8750 1.0800 2.0450 1.2050 ;
	    RECT 1.8750 0.8700 2.3650 1.0800 ;
	    RECT 2.1950 0.5300 2.3650 0.8700 ;
	    RECT 2.5400 0.7450 2.7100 1.9200 ;
	    RECT 3.7050 1.6550 3.8750 1.9200 ;
	    RECT 4.0450 2.1200 4.2150 2.3700 ;
	    RECT 4.0450 1.9050 4.5550 2.1200 ;
	    RECT 4.2000 1.7200 4.5550 1.9050 ;
	    RECT 3.7050 1.2450 4.0300 1.6550 ;
	    RECT 2.9900 0.7650 4.0300 0.9350 ;
	    RECT 3.4100 0.5300 3.6900 0.5950 ;
	    RECT 2.1950 0.2650 3.6900 0.5300 ;
	    RECT 3.8600 0.5300 4.0300 0.7650 ;
	    RECT 4.2000 0.7450 4.3700 1.7200 ;
	    RECT 4.7250 1.5050 4.8950 2.3700 ;
	    RECT 5.1250 1.8050 5.5400 2.1450 ;
	    RECT 4.5400 1.3150 4.8950 1.5050 ;
	    RECT 4.5400 1.3050 4.8900 1.3150 ;
	    RECT 4.5400 1.3000 4.8800 1.3050 ;
	    RECT 4.5400 1.2950 4.8650 1.3000 ;
	    RECT 4.5400 0.5300 4.7100 1.2950 ;
	    RECT 3.8600 0.3200 4.7100 0.5300 ;
	    RECT 5.3000 0.5200 5.5400 1.8050 ;
	    RECT 5.7150 0.7450 5.8850 2.6300 ;
	    RECT 6.0750 1.1150 6.2450 2.8450 ;
	    RECT 9.4150 2.6300 9.7350 3.0800 ;
	    RECT 6.4150 2.0200 6.8300 2.5550 ;
	    RECT 7.1650 2.4200 9.7350 2.6300 ;
	    RECT 6.4150 1.8050 6.9950 2.0200 ;
	    RECT 6.4300 1.2450 6.6550 1.5950 ;
	    RECT 6.0750 0.9000 6.3150 1.1150 ;
	    RECT 6.4850 0.9900 6.6550 1.2450 ;
	    RECT 6.1100 0.8300 6.3150 0.9000 ;
	    RECT 6.1100 0.7550 6.4000 0.8300 ;
	    RECT 5.7150 0.6450 5.9350 0.7450 ;
	    RECT 5.7150 0.3150 5.9800 0.6450 ;
	    RECT 6.1500 0.4000 6.4000 0.7550 ;
	    RECT 6.8250 0.5300 6.9950 1.8050 ;
	    RECT 7.1650 0.7450 7.3350 2.4200 ;
	    RECT 9.1900 2.3450 9.7350 2.4200 ;
	    RECT 8.4550 1.8700 9.3950 2.1300 ;
	    RECT 8.0450 1.1800 8.2550 1.5950 ;
	    RECT 8.0450 0.9150 8.2500 1.1800 ;
	    RECT 9.2250 1.1300 9.3950 1.8700 ;
	    RECT 8.5350 0.9400 9.3950 1.1300 ;
	    RECT 8.4950 0.9200 9.3950 0.9400 ;
	    RECT 7.7050 0.5300 8.1700 0.5800 ;
	    RECT 6.8250 0.3200 8.1700 0.5300 ;
	    RECT 8.4950 0.3700 8.7850 0.9200 ;
	    RECT 9.5650 0.7300 9.7350 2.3450 ;
	    RECT 9.4150 0.3200 9.7350 0.7300 ;
         LAYER met1 ;
	    RECT 4.3250 2.0000 4.6150 2.0550 ;
	    RECT 6.6250 2.0000 6.9150 2.0550 ;
	    RECT 4.3250 1.8250 6.9150 2.0000 ;
	    RECT 4.3250 1.7700 4.6150 1.8250 ;
	    RECT 6.6250 1.7700 6.9150 1.8250 ;
	    RECT 5.2450 1.1900 5.5350 1.2050 ;
	    RECT 6.4850 1.1900 6.9150 1.2050 ;
	    RECT 5.2450 1.1500 6.9150 1.1900 ;
	    RECT 8.0050 1.1500 8.2950 1.2050 ;
	    RECT 5.2450 0.9750 8.2950 1.1500 ;
	    RECT 5.2450 0.9600 6.9150 0.9750 ;
	    RECT 5.2450 0.9200 5.5350 0.9600 ;
	    RECT 6.4850 0.9200 6.9150 0.9600 ;
	    RECT 8.0050 0.9200 8.2950 0.9750 ;
	    RECT 5.7050 0.7250 5.9950 0.7800 ;
	    RECT 8.4650 0.7250 8.7550 0.7800 ;
	    RECT 5.7050 0.5500 8.7550 0.7250 ;
	    RECT 5.7050 0.4950 5.9950 0.5500 ;
	    RECT 8.4650 0.4950 8.7550 0.5500 ;
   END
END efs8hd_xor3_4
MACRO efs8hd_clkbuf_1
   CLASS CORE ;
   FOREIGN efs8hd_clkbuf_1 ;
   ORIGIN -0.0000 -0.0000 ;
   SIZE 1.3800 BY 3.4000 ;
   PIN A
      PORT
         LAYER li1 ;
	    RECT 0.9450 1.2300 1.2750 1.6900 ;
      END
   END A
   PIN X
      PORT
         LAYER li1 ;
	    RECT 0.0850 1.9500 0.3550 3.0800 ;
	    RECT 0.0850 0.9500 0.2550 1.9500 ;
	    RECT 0.0850 0.3150 0.3450 0.9500 ;
      END
   END X
   PIN vgnd
      PORT
         LAYER li1 ;
	    RECT 0.5250 0.0850 0.8550 0.5800 ;
	    RECT 0.0000 -0.0850 1.3800 0.0850 ;
         LAYER met1 ;
	    RECT 0.0000 -0.3000 1.3800 0.3000 ;
      END
   END vgnd
   PIN vpwr
      PORT
         LAYER li1 ;
	    RECT 0.0000 3.3150 1.3800 3.4850 ;
	    RECT 0.5250 2.3400 0.8550 3.3150 ;
         LAYER met1 ;
	    RECT 0.0000 3.1000 1.3800 3.7000 ;
      END
   END vpwr
   OBS
         LAYER li1 ;
	    RECT 1.0350 2.1300 1.2050 3.0800 ;
	    RECT 0.5400 1.9150 1.2050 2.1300 ;
	    RECT 0.5400 1.7350 0.7100 1.9150 ;
	    RECT 0.4250 1.3250 0.7100 1.7350 ;
	    RECT 0.5400 1.0050 0.7100 1.3250 ;
	    RECT 0.5400 0.7900 1.2050 1.0050 ;
	    RECT 1.0350 0.3150 1.2050 0.7900 ;
   END
END efs8hd_clkbuf_1
END LIBRARY
