// Copyright 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

(* blackbox *)
module sky130_fd_sc_hd__dfrbp_1  (output QN, input D, input CLK, output Q, input RESETB); endmodule
(* blackbox *)
module sky130_fd_sc_hd__inv_4 (input A, output Y); endmodule
(* blackbox *)
module sky130_fd_sc_hd__buf_1(input A, output X); endmodule
(* blackbox *)
module sky130_fd_sc_hd__clkbuf_1(input A, output X); endmodule
(* blackbox *)
module sky130_fd_sc_hd__clkbuf_2(input A, output X); endmodule
(* blackbox *)
module sky130_fd_sc_hd__clkinv_1(input A, output Y); endmodule
(* blackbox *)
module sky130_fd_sc_hd__clkinv_2(input A, output Y); endmodule
(* blackbox *)
module sky130_fd_sc_hd__clkinv_4(input A, output Y); endmodule
(* blackbox *)
module sky130_fd_sc_hd__clkinv_8(input A, output Y); endmodule
(* blackbox *)
module sky130_fd_sc_hd__conb_1(output HI, output LO); endmodule
(* blackbox *)
module sky130_fd_sc_hd__dfbbp_1(input CLK, input D, output Q, output QN, input RESETB, input SETB); endmodule
(* blackbox *)
module sky130_fd_sc_hd__einvn_4(input A, input TEB, output Z); endmodule
(* blackbox *)
module sky130_fd_sc_hd__einvn_8(input A, input TEB, output Z); endmodule
(* blackbox *)
module sky130_fd_sc_hd__einvp_1(input A, input TE, output Z); endmodule
(* blackbox *)
module sky130_fd_sc_hd__einvp_2(input A, input TE, output Z); endmodule
(* blackbox *)
module sky130_fd_sc_hd__or2_2(input A, B, output X); endmodule
