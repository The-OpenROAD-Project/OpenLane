(* blackbox *)
module scs8hd_inv_1 (input A, output Y); endmodule
(* blackbox *)
module scs8hd_inv_2 (input A, output Y); endmodule
(* blackbox *)
module scs8hd_inv_4 (input A, output Y); endmodule
(* blackbox *)
module scs8hd_buf_1(input A, output X); endmodule
(* blackbox *)
module scs8hd_buf_2(input A, output X); endmodule
(* blackbox *)
module scs8hd_buf_4(input A, output X); endmodule
(* blackbox *)
module scs8hd_or2_1(input A, input B, output X); endmodule
(* blackbox *)
module scs8hd_mux2_1(input A0, input A1, input S, output X); endmodule
(* blackbox *)
module scs8hd_dfrtp_1(input CLK, input D, input RESETB, output Q); endmodule
(* blackbox *)
module scs8hd_dfrbp_1(input CLK, input D, input RESETB, output Q, output QN); endmodule
(* blackbox *)
module iopad(input en, input inpad, output outpad, output pad); endmodule



