magic
tech sky130A
magscale 1 2
timestamp 1636140361
<< checkpaint >>
rect -1296 -1277 3932 2731
<< nwell >>
rect -36 679 2672 1471
<< locali >>
rect 0 1397 2636 1431
rect 64 674 98 740
rect 1263 690 1297 724
rect 0 -17 2636 17
use sky130_sram_1kbyte_1rw1r_32x256_8_pinv_15  sky130_sram_1kbyte_1rw1r_32x256_8_pinv_15_0
timestamp 1636140361
transform 1 0 0 0 1 0
box -36 -17 2672 1471
<< labels >>
rlabel locali s 1280 707 1280 707 4 Z
port 1 nsew
rlabel locali s 81 707 81 707 4 A
port 2 nsew
rlabel locali s 1318 0 1318 0 4 gnd
port 3 nsew
rlabel locali s 1318 1414 1318 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2636 1414
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_END 358828
string GDS_START 357996
<< end >>
