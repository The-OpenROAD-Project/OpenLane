magic
tech sky130A
magscale 1 2
timestamp 1636140361
<< checkpaint >>
rect -1296 -1277 2438 2731
<< nwell >>
rect -36 679 1178 1471
<< locali >>
rect 0 1397 1142 1431
rect 64 636 98 702
rect 179 671 449 705
rect 805 690 965 724
rect 1063 690 1097 724
rect 547 687 581 688
rect 179 669 213 671
rect 547 653 707 687
rect 805 670 839 690
rect 0 -17 1142 17
use pinv_19  pinv_19_0
timestamp 1636140361
transform 1 0 884 0 1 0
box -36 -17 294 1471
use pinv_18  pinv_18_0
timestamp 1636140361
transform 1 0 626 0 1 0
box -36 -17 294 1471
use pinv_12  pinv_12_0
timestamp 1636140361
transform 1 0 368 0 1 0
box -36 -17 294 1471
use pinv_6  pinv_6_0
timestamp 1636140361
transform 1 0 0 0 1 0
box -36 -17 404 1471
<< labels >>
rlabel locali s 1080 707 1080 707 4 Z
port 2 nsew
rlabel locali s 81 669 81 669 4 A
port 1 nsew
rlabel locali s 571 1414 571 1414 4 vdd
port 3 nsew
rlabel locali s 571 0 571 0 4 gnd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1142 1414
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_END 4886532
string GDS_START 4885022
<< end >>
