magic
tech sky130A
magscale 1 2
timestamp 1636140361
<< checkpaint >>
rect -1260 -1260 1261 1261
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_END 4737978
string GDS_START 4737654
<< end >>
