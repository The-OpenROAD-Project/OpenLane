VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO sram_1rw1r_32_256_8_s8
  CLASS BLOCK ;
  FOREIGN sram_1rw1r_32_256_8_s8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 390.820 BY 574.890 ;
  SYMMETRY X Y R90 ;
  PIN din0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.745 5.440 80.075 9.700 ;
    END
  END din0[0]


  PIN din0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.575 5.440 85.905 9.700 ;
    END
  END din0[1]


  PIN din0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.405 5.440 91.735 9.700 ;
    END
  END din0[2]


  PIN din0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.235 5.440 97.565 9.700 ;
    END
  END din0[3]


  PIN din0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.065 5.440 103.395 9.700 ;
    END
  END din0[4]


  PIN din0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.895 5.440 109.225 9.700 ;
    END
  END din0[5]


  PIN din0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 114.725 5.440 115.055 9.700 ;
    END
  END din0[6]


  PIN din0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 120.555 5.440 120.885 9.700 ;
    END
  END din0[7]


  PIN din0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.385 5.440 126.715 9.700 ;
    END
  END din0[8]


  PIN din0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.215 5.440 132.545 9.700 ;
    END
  END din0[9]


  PIN din0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.045 5.440 138.375 9.700 ;
    END
  END din0[10]


  PIN din0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.875 5.440 144.205 9.700 ;
    END
  END din0[11]


  PIN din0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.705 5.440 150.035 9.700 ;
    END
  END din0[12]


  PIN din0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.535 5.440 155.865 9.700 ;
    END
  END din0[13]


  PIN din0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 161.365 5.440 161.695 9.700 ;
    END
  END din0[14]


  PIN din0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 167.195 5.440 167.525 9.700 ;
    END
  END din0[15]


  PIN din0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.025 5.440 173.355 9.700 ;
    END
  END din0[16]


  PIN din0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.855 5.440 179.185 9.700 ;
    END
  END din0[17]


  PIN din0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 184.685 5.440 185.015 9.700 ;
    END
  END din0[18]


  PIN din0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.515 5.440 190.845 9.700 ;
    END
  END din0[19]


  PIN din0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 196.345 5.440 196.675 9.700 ;
    END
  END din0[20]


  PIN din0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.175 5.440 202.505 9.700 ;
    END
  END din0[21]


  PIN din0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.005 5.440 208.335 9.700 ;
    END
  END din0[22]


  PIN din0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 213.835 5.440 214.165 9.700 ;
    END
  END din0[23]


  PIN din0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 219.665 5.440 219.995 9.700 ;
    END
  END din0[24]


  PIN din0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 225.495 5.440 225.825 9.700 ;
    END
  END din0[25]


  PIN din0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.325 5.440 231.655 9.700 ;
    END
  END din0[26]


  PIN din0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 237.155 5.440 237.485 9.700 ;
    END
  END din0[27]


  PIN din0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.985 5.440 243.315 9.700 ;
    END
  END din0[28]


  PIN din0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 248.815 5.440 249.145 9.700 ;
    END
  END din0[29]


  PIN din0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.645 5.440 254.975 9.700 ;
    END
  END din0[30]


  PIN din0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 260.475 5.440 260.805 9.700 ;
    END
  END din0[31]


  PIN addr0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.655 5.440 72.985 9.700 ;
    END
  END addr0[0]


  PIN addr0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.140 402.865 9.700 403.125 ;
    END
  END addr0[1]


  PIN addr0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.140 411.385 9.700 411.645 ;
    END
  END addr0[2]


  PIN addr0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.140 417.005 9.700 417.265 ;
    END
  END addr0[3]


  PIN addr0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.140 425.525 9.700 425.785 ;
    END
  END addr0[4]


  PIN addr0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.140 431.145 9.700 431.405 ;
    END
  END addr0[5]


  PIN addr0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.140 439.665 9.700 439.925 ;
    END
  END addr0[6]


  PIN addr0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.140 445.285 9.700 445.545 ;
    END
  END addr0[7]


  PIN addr1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.120 457.375 386.680 457.635 ;
    END
  END addr1[0]


  PIN addr1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.120 115.740 386.680 116.000 ;
    END
  END addr1[1]


  PIN addr1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.120 107.220 386.680 107.480 ;
    END
  END addr1[2]


  PIN addr1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.120 101.600 386.680 101.860 ;
    END
  END addr1[3]


  PIN addr1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.120 93.080 386.680 93.340 ;
    END
  END addr1[4]


  PIN addr1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.120 87.460 386.680 87.720 ;
    END
  END addr1[5]


  PIN addr1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.120 78.940 386.680 79.200 ;
    END
  END addr1[6]


  PIN addr1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.120 73.320 386.680 73.580 ;
    END
  END addr1[7]


  PIN csb0
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.140 54.690 9.700 54.950 ;
    END
  END csb0


  PIN csb1
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.120 467.530 386.680 467.790 ;
    END
  END csb1


  PIN web0
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.140 63.210 9.700 63.470 ;
    END
  END web0


  PIN clk0
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.535 5.440 23.675 9.700 ;
    END
  END clk0


  PIN clk1
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 346.945 565.190 347.085 569.450 ;
    END
  END clk1


  PIN wmask0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.300 5.440 67.630 9.700 ;
    END
  END wmask0[0]


  PIN wmask0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.750 5.440 62.080 9.700 ;
    END
  END wmask0[1]


  PIN wmask0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.305 5.440 55.635 9.700 ;
    END
  END wmask0[2]


  PIN wmask0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.885 5.440 46.215 9.700 ;
    END
  END wmask0[3]


  PIN dout0[0]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 85.820 5.440 86.035 9.700 ;
    END
  END dout0[0]


  PIN dout0[1]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 92.060 5.440 92.275 9.700 ;
    END
  END dout0[1]


  PIN dout0[2]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 98.300 5.440 98.515 9.700 ;
    END
  END dout0[2]


  PIN dout0[3]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 105.780 5.440 105.920 9.700 ;
    END
  END dout0[3]


  PIN dout0[4]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 112.020 5.440 112.160 9.700 ;
    END
  END dout0[4]


  PIN dout0[5]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 117.020 5.440 117.235 9.700 ;
    END
  END dout0[5]


  PIN dout0[6]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 123.260 5.440 123.475 9.700 ;
    END
  END dout0[6]


  PIN dout0[7]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 130.740 5.440 130.880 9.700 ;
    END
  END dout0[7]


  PIN dout0[8]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 136.980 5.440 137.120 9.700 ;
    END
  END dout0[8]


  PIN dout0[9]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 141.980 5.440 142.195 9.700 ;
    END
  END dout0[9]


  PIN dout0[10]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 148.220 5.440 148.435 9.700 ;
    END
  END dout0[10]


  PIN dout0[11]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 155.700 5.440 155.840 9.700 ;
    END
  END dout0[11]


  PIN dout0[12]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 161.940 5.440 162.080 9.700 ;
    END
  END dout0[12]


  PIN dout0[13]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 166.940 5.440 167.155 9.700 ;
    END
  END dout0[13]


  PIN dout0[14]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 173.180 5.440 173.395 9.700 ;
    END
  END dout0[14]


  PIN dout0[15]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 180.660 5.440 180.800 9.700 ;
    END
  END dout0[15]


  PIN dout0[16]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 186.900 5.440 187.040 9.700 ;
    END
  END dout0[16]


  PIN dout0[17]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 191.900 5.440 192.115 9.700 ;
    END
  END dout0[17]


  PIN dout0[18]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 198.140 5.440 198.355 9.700 ;
    END
  END dout0[18]


  PIN dout0[19]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 205.620 5.440 205.760 9.700 ;
    END
  END dout0[19]


  PIN dout0[20]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 211.860 5.440 212.000 9.700 ;
    END
  END dout0[20]


  PIN dout0[21]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 216.860 5.440 217.075 9.700 ;
    END
  END dout0[21]


  PIN dout0[22]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 223.100 5.440 223.315 9.700 ;
    END
  END dout0[22]


  PIN dout0[23]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 230.580 5.440 230.720 9.700 ;
    END
  END dout0[23]


  PIN dout0[24]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 236.820 5.440 236.960 9.700 ;
    END
  END dout0[24]


  PIN dout0[25]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 241.820 5.440 242.035 9.700 ;
    END
  END dout0[25]


  PIN dout0[26]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 248.060 5.440 248.275 9.700 ;
    END
  END dout0[26]


  PIN dout0[27]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 255.540 5.440 255.680 9.700 ;
    END
  END dout0[27]


  PIN dout0[28]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 261.780 5.440 261.920 9.700 ;
    END
  END dout0[28]


  PIN dout0[29]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 266.780 5.440 266.995 9.700 ;
    END
  END dout0[29]


  PIN dout0[30]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 273.020 5.440 273.235 9.700 ;
    END
  END dout0[30]


  PIN dout0[31]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 280.500 5.440 280.640 9.700 ;
    END
  END dout0[31]


  PIN dout1[0]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 85.820 565.190 85.960 569.450 ;
    END
  END dout1[0]


  PIN dout1[1]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 92.060 565.190 92.200 569.450 ;
    END
  END dout1[1]


  PIN dout1[2]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 98.300 565.190 98.440 569.450 ;
    END
  END dout1[2]


  PIN dout1[3]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 105.780 565.190 105.920 569.450 ;
    END
  END dout1[3]


  PIN dout1[4]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 112.020 565.190 112.160 569.450 ;
    END
  END dout1[4]


  PIN dout1[5]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 117.020 565.190 117.160 569.450 ;
    END
  END dout1[5]


  PIN dout1[6]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 123.260 565.190 123.400 569.450 ;
    END
  END dout1[6]


  PIN dout1[7]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 130.740 565.190 130.880 569.450 ;
    END
  END dout1[7]


  PIN dout1[8]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 136.980 565.190 137.120 569.450 ;
    END
  END dout1[8]


  PIN dout1[9]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 141.980 565.190 142.120 569.450 ;
    END
  END dout1[9]


  PIN dout1[10]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 148.220 565.190 148.360 569.450 ;
    END
  END dout1[10]


  PIN dout1[11]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 155.700 565.190 155.840 569.450 ;
    END
  END dout1[11]


  PIN dout1[12]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 161.940 565.190 162.080 569.450 ;
    END
  END dout1[12]


  PIN dout1[13]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 166.940 565.190 167.080 569.450 ;
    END
  END dout1[13]


  PIN dout1[14]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 173.180 565.190 173.320 569.450 ;
    END
  END dout1[14]


  PIN dout1[15]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 180.660 565.190 180.800 569.450 ;
    END
  END dout1[15]


  PIN dout1[16]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 186.900 565.190 187.040 569.450 ;
    END
  END dout1[16]


  PIN dout1[17]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 191.900 565.190 192.040 569.450 ;
    END
  END dout1[17]


  PIN dout1[18]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 198.140 565.190 198.280 569.450 ;
    END
  END dout1[18]


  PIN dout1[19]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 205.620 565.190 205.760 569.450 ;
    END
  END dout1[19]


  PIN dout1[20]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 211.860 565.190 212.000 569.450 ;
    END
  END dout1[20]


  PIN dout1[21]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 216.860 565.190 217.000 569.450 ;
    END
  END dout1[21]


  PIN dout1[22]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 223.100 565.190 223.240 569.450 ;
    END
  END dout1[22]


  PIN dout1[23]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 230.580 565.190 230.720 569.450 ;
    END
  END dout1[23]


  PIN dout1[24]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 236.820 565.190 236.960 569.450 ;
    END
  END dout1[24]


  PIN dout1[25]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 241.820 565.190 241.960 569.450 ;
    END
  END dout1[25]


  PIN dout1[26]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 248.060 565.190 248.200 569.450 ;
    END
  END dout1[26]


  PIN dout1[27]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 255.540 565.190 255.680 569.450 ;
    END
  END dout1[27]


  PIN dout1[28]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 261.780 565.190 261.920 569.450 ;
    END
  END dout1[28]


  PIN dout1[29]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 266.780 565.190 266.920 569.450 ;
    END
  END dout1[29]


  PIN dout1[30]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 273.020 565.190 273.160 569.450 ;
    END
  END dout1[30]


  PIN dout1[31]
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 280.500 565.190 280.640 569.450 ;
    END
  END dout1[31]


  OBS
     LAYER li1 ;
       RECT 10.000 10.000 380.82 564.89 ;
     LAYER met1 ;
       RECT 10.000 10.000 380.82 564.89 ;
     LAYER met2 ;
       RECT 10.000 10.000 380.82 564.89 ;
     LAYER met3 ;
       RECT 10.000 10.000 380.82 564.89 ;
     LAYER met4 ;
       RECT 10.000 10.000 380.82 564.89 ;
     LAYER met5 ;
       RECT 10.000 10.000 380.82 564.89 ;
  END
END sram_1rw1r_32_256_8_s8
