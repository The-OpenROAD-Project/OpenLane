magic
tech sky130A
magscale 1 2
timestamp 1636140361
<< checkpaint >>
rect -1260 -1260 68594 68572
<< locali >>
rect 60352 66122 60386 66138
rect 60352 66072 60386 66088
rect 59953 65415 59987 65431
rect 61039 65419 61073 65453
rect 59953 65365 59987 65381
rect 60352 64708 60386 64724
rect 60352 64658 60386 64674
rect 59953 64001 59987 64017
rect 59953 63951 59987 63967
rect 60352 63294 60386 63310
rect 60352 63244 60386 63260
rect 55077 60873 55111 60889
rect 55111 60839 55257 60873
rect 55077 60823 55111 60839
rect 12139 60633 12173 60649
rect 11993 60599 12139 60633
rect 12139 60583 12173 60599
rect 55077 60633 55111 60649
rect 55111 60599 55257 60633
rect 55077 60583 55111 60599
rect 12139 60083 12173 60099
rect 11993 60049 12139 60083
rect 12139 60033 12173 60049
rect 55077 60083 55111 60099
rect 55111 60049 55257 60083
rect 55077 60033 55111 60049
rect 12139 59843 12173 59859
rect 11993 59809 12139 59843
rect 12139 59793 12173 59809
rect 55077 59843 55111 59859
rect 55111 59809 55257 59843
rect 55077 59793 55111 59809
rect 12139 59293 12173 59309
rect 11993 59259 12139 59293
rect 12139 59243 12173 59259
rect 55077 59293 55111 59309
rect 55111 59259 55257 59293
rect 55077 59243 55111 59259
rect 12139 59053 12173 59069
rect 11993 59019 12139 59053
rect 12139 59003 12173 59019
rect 55077 59053 55111 59069
rect 55111 59019 55257 59053
rect 55077 59003 55111 59019
rect 12139 58503 12173 58519
rect 11993 58469 12139 58503
rect 12139 58453 12173 58469
rect 55077 58503 55111 58519
rect 55111 58469 55257 58503
rect 55077 58453 55111 58469
rect 12139 58263 12173 58279
rect 11993 58229 12139 58263
rect 12139 58213 12173 58229
rect 55077 58263 55111 58279
rect 55111 58229 55257 58263
rect 55077 58213 55111 58229
rect 12139 57713 12173 57729
rect 11993 57679 12139 57713
rect 12139 57663 12173 57679
rect 55077 57713 55111 57729
rect 55111 57679 55257 57713
rect 55077 57663 55111 57679
rect 12139 57473 12173 57489
rect 11993 57439 12139 57473
rect 12139 57423 12173 57439
rect 55077 57473 55111 57489
rect 55111 57439 55257 57473
rect 55077 57423 55111 57439
rect 12139 56923 12173 56939
rect 11993 56889 12139 56923
rect 12139 56873 12173 56889
rect 55077 56923 55111 56939
rect 55111 56889 55257 56923
rect 55077 56873 55111 56889
rect 12139 56683 12173 56699
rect 11993 56649 12139 56683
rect 12139 56633 12173 56649
rect 55077 56683 55111 56699
rect 55111 56649 55257 56683
rect 55077 56633 55111 56649
rect 12139 56133 12173 56149
rect 11993 56099 12139 56133
rect 12139 56083 12173 56099
rect 55077 56133 55111 56149
rect 55111 56099 55257 56133
rect 55077 56083 55111 56099
rect 12139 55893 12173 55909
rect 11993 55859 12139 55893
rect 12139 55843 12173 55859
rect 55077 55893 55111 55909
rect 55111 55859 55257 55893
rect 55077 55843 55111 55859
rect 12139 55343 12173 55359
rect 11993 55309 12139 55343
rect 12139 55293 12173 55309
rect 55077 55343 55111 55359
rect 55111 55309 55257 55343
rect 55077 55293 55111 55309
rect 12139 55103 12173 55119
rect 11993 55069 12139 55103
rect 12139 55053 12173 55069
rect 55077 55103 55111 55119
rect 55111 55069 55257 55103
rect 55077 55053 55111 55069
rect 12139 54553 12173 54569
rect 11993 54519 12139 54553
rect 12139 54503 12173 54519
rect 55077 54553 55111 54569
rect 55111 54519 55257 54553
rect 55077 54503 55111 54519
rect 12139 54313 12173 54329
rect 11993 54279 12139 54313
rect 12139 54263 12173 54279
rect 55077 54313 55111 54329
rect 55111 54279 55257 54313
rect 55077 54263 55111 54279
rect 12139 53763 12173 53779
rect 11993 53729 12139 53763
rect 12139 53713 12173 53729
rect 55077 53763 55111 53779
rect 55111 53729 55257 53763
rect 55077 53713 55111 53729
rect 12139 53523 12173 53539
rect 11993 53489 12139 53523
rect 12139 53473 12173 53489
rect 55077 53523 55111 53539
rect 55111 53489 55257 53523
rect 55077 53473 55111 53489
rect 12139 52973 12173 52989
rect 11993 52939 12139 52973
rect 12139 52923 12173 52939
rect 55077 52973 55111 52989
rect 55111 52939 55257 52973
rect 55077 52923 55111 52939
rect 12139 52733 12173 52749
rect 11993 52699 12139 52733
rect 12139 52683 12173 52699
rect 55077 52733 55111 52749
rect 55111 52699 55257 52733
rect 55077 52683 55111 52699
rect 12139 52183 12173 52199
rect 11993 52149 12139 52183
rect 12139 52133 12173 52149
rect 55077 52183 55111 52199
rect 55111 52149 55257 52183
rect 55077 52133 55111 52149
rect 12139 51943 12173 51959
rect 11993 51909 12139 51943
rect 12139 51893 12173 51909
rect 55077 51943 55111 51959
rect 55111 51909 55257 51943
rect 55077 51893 55111 51909
rect 12139 51393 12173 51409
rect 11993 51359 12139 51393
rect 12139 51343 12173 51359
rect 55077 51393 55111 51409
rect 55111 51359 55257 51393
rect 55077 51343 55111 51359
rect 12139 51153 12173 51169
rect 11993 51119 12139 51153
rect 12139 51103 12173 51119
rect 55077 51153 55111 51169
rect 55111 51119 55257 51153
rect 55077 51103 55111 51119
rect 12139 50603 12173 50619
rect 11993 50569 12139 50603
rect 12139 50553 12173 50569
rect 55077 50603 55111 50619
rect 55111 50569 55257 50603
rect 55077 50553 55111 50569
rect 12139 50363 12173 50379
rect 11993 50329 12139 50363
rect 12139 50313 12173 50329
rect 55077 50363 55111 50379
rect 55111 50329 55257 50363
rect 55077 50313 55111 50329
rect 12139 49813 12173 49829
rect 11993 49779 12139 49813
rect 12139 49763 12173 49779
rect 55077 49813 55111 49829
rect 55111 49779 55257 49813
rect 55077 49763 55111 49779
rect 12139 49573 12173 49589
rect 11993 49539 12139 49573
rect 12139 49523 12173 49539
rect 55077 49573 55111 49589
rect 55111 49539 55257 49573
rect 55077 49523 55111 49539
rect 12139 49023 12173 49039
rect 11993 48989 12139 49023
rect 12139 48973 12173 48989
rect 55077 49023 55111 49039
rect 55111 48989 55257 49023
rect 55077 48973 55111 48989
rect 12139 48783 12173 48799
rect 11993 48749 12139 48783
rect 12139 48733 12173 48749
rect 55077 48783 55111 48799
rect 55111 48749 55257 48783
rect 55077 48733 55111 48749
rect 12139 48233 12173 48249
rect 11993 48199 12139 48233
rect 12139 48183 12173 48199
rect 55077 48233 55111 48249
rect 55111 48199 55257 48233
rect 55077 48183 55111 48199
rect 12139 47993 12173 48009
rect 11993 47959 12139 47993
rect 12139 47943 12173 47959
rect 55077 47993 55111 48009
rect 55111 47959 55257 47993
rect 55077 47943 55111 47959
rect 12139 47443 12173 47459
rect 11993 47409 12139 47443
rect 12139 47393 12173 47409
rect 55077 47443 55111 47459
rect 55111 47409 55257 47443
rect 55077 47393 55111 47409
rect 12139 47203 12173 47219
rect 11993 47169 12139 47203
rect 12139 47153 12173 47169
rect 55077 47203 55111 47219
rect 55111 47169 55257 47203
rect 55077 47153 55111 47169
rect 12139 46653 12173 46669
rect 11993 46619 12139 46653
rect 12139 46603 12173 46619
rect 55077 46653 55111 46669
rect 55111 46619 55257 46653
rect 55077 46603 55111 46619
rect 12139 46413 12173 46429
rect 11993 46379 12139 46413
rect 12139 46363 12173 46379
rect 55077 46413 55111 46429
rect 55111 46379 55257 46413
rect 55077 46363 55111 46379
rect 12139 45863 12173 45879
rect 11993 45829 12139 45863
rect 12139 45813 12173 45829
rect 55077 45863 55111 45879
rect 55111 45829 55257 45863
rect 55077 45813 55111 45829
rect 12139 45623 12173 45639
rect 11993 45589 12139 45623
rect 12139 45573 12173 45589
rect 55077 45623 55111 45639
rect 55111 45589 55257 45623
rect 55077 45573 55111 45589
rect 12139 45073 12173 45089
rect 11993 45039 12139 45073
rect 12139 45023 12173 45039
rect 55077 45073 55111 45089
rect 55111 45039 55257 45073
rect 55077 45023 55111 45039
rect 12139 44833 12173 44849
rect 11993 44799 12139 44833
rect 12139 44783 12173 44799
rect 55077 44833 55111 44849
rect 55111 44799 55257 44833
rect 55077 44783 55111 44799
rect 12139 44283 12173 44299
rect 11993 44249 12139 44283
rect 12139 44233 12173 44249
rect 55077 44283 55111 44299
rect 55111 44249 55257 44283
rect 55077 44233 55111 44249
rect 12139 44043 12173 44059
rect 11993 44009 12139 44043
rect 12139 43993 12173 44009
rect 55077 44043 55111 44059
rect 55111 44009 55257 44043
rect 55077 43993 55111 44009
rect 12139 43493 12173 43509
rect 11993 43459 12139 43493
rect 12139 43443 12173 43459
rect 55077 43493 55111 43509
rect 55111 43459 55257 43493
rect 55077 43443 55111 43459
rect 12139 43253 12173 43269
rect 11993 43219 12139 43253
rect 12139 43203 12173 43219
rect 55077 43253 55111 43269
rect 55111 43219 55257 43253
rect 55077 43203 55111 43219
rect 12139 42703 12173 42719
rect 11993 42669 12139 42703
rect 12139 42653 12173 42669
rect 55077 42703 55111 42719
rect 55111 42669 55257 42703
rect 55077 42653 55111 42669
rect 12139 42463 12173 42479
rect 11993 42429 12139 42463
rect 12139 42413 12173 42429
rect 55077 42463 55111 42479
rect 55111 42429 55257 42463
rect 55077 42413 55111 42429
rect 12139 41913 12173 41929
rect 11993 41879 12139 41913
rect 12139 41863 12173 41879
rect 55077 41913 55111 41929
rect 55111 41879 55257 41913
rect 55077 41863 55111 41879
rect 12139 41673 12173 41689
rect 11993 41639 12139 41673
rect 12139 41623 12173 41639
rect 55077 41673 55111 41689
rect 55111 41639 55257 41673
rect 55077 41623 55111 41639
rect 12139 41123 12173 41139
rect 11993 41089 12139 41123
rect 12139 41073 12173 41089
rect 55077 41123 55111 41139
rect 55111 41089 55257 41123
rect 55077 41073 55111 41089
rect 12139 40883 12173 40899
rect 11993 40849 12139 40883
rect 12139 40833 12173 40849
rect 55077 40883 55111 40899
rect 55111 40849 55257 40883
rect 55077 40833 55111 40849
rect 12139 40333 12173 40349
rect 11993 40299 12139 40333
rect 12139 40283 12173 40299
rect 55077 40333 55111 40349
rect 55111 40299 55257 40333
rect 55077 40283 55111 40299
rect 12139 40093 12173 40109
rect 11993 40059 12139 40093
rect 12139 40043 12173 40059
rect 55077 40093 55111 40109
rect 55111 40059 55257 40093
rect 55077 40043 55111 40059
rect 12139 39543 12173 39559
rect 11993 39509 12139 39543
rect 12139 39493 12173 39509
rect 55077 39543 55111 39559
rect 55111 39509 55257 39543
rect 55077 39493 55111 39509
rect 12139 39303 12173 39319
rect 11993 39269 12139 39303
rect 12139 39253 12173 39269
rect 55077 39303 55111 39319
rect 55111 39269 55257 39303
rect 55077 39253 55111 39269
rect 12139 38753 12173 38769
rect 11993 38719 12139 38753
rect 12139 38703 12173 38719
rect 55077 38753 55111 38769
rect 55111 38719 55257 38753
rect 55077 38703 55111 38719
rect 12139 38513 12173 38529
rect 11993 38479 12139 38513
rect 12139 38463 12173 38479
rect 55077 38513 55111 38529
rect 55111 38479 55257 38513
rect 55077 38463 55111 38479
rect 12139 37963 12173 37979
rect 11993 37929 12139 37963
rect 12139 37913 12173 37929
rect 55077 37963 55111 37979
rect 55111 37929 55257 37963
rect 55077 37913 55111 37929
rect 12139 37723 12173 37739
rect 11993 37689 12139 37723
rect 12139 37673 12173 37689
rect 55077 37723 55111 37739
rect 55111 37689 55257 37723
rect 55077 37673 55111 37689
rect 12139 37173 12173 37189
rect 11993 37139 12139 37173
rect 12139 37123 12173 37139
rect 55077 37173 55111 37189
rect 55111 37139 55257 37173
rect 55077 37123 55111 37139
rect 12139 36933 12173 36949
rect 11993 36899 12139 36933
rect 12139 36883 12173 36899
rect 55077 36933 55111 36949
rect 55111 36899 55257 36933
rect 55077 36883 55111 36899
rect 12139 36383 12173 36399
rect 11993 36349 12139 36383
rect 12139 36333 12173 36349
rect 55077 36383 55111 36399
rect 55111 36349 55257 36383
rect 55077 36333 55111 36349
rect 12139 36143 12173 36159
rect 11993 36109 12139 36143
rect 12139 36093 12173 36109
rect 55077 36143 55111 36159
rect 55111 36109 55257 36143
rect 55077 36093 55111 36109
rect 12139 35593 12173 35609
rect 11993 35559 12139 35593
rect 12139 35543 12173 35559
rect 55077 35593 55111 35609
rect 55111 35559 55257 35593
rect 55077 35543 55111 35559
rect 12139 35353 12173 35369
rect 11993 35319 12139 35353
rect 12139 35303 12173 35319
rect 55077 35353 55111 35369
rect 55111 35319 55257 35353
rect 55077 35303 55111 35319
rect 12139 34803 12173 34819
rect 11993 34769 12139 34803
rect 12139 34753 12173 34769
rect 55077 34803 55111 34819
rect 55111 34769 55257 34803
rect 55077 34753 55111 34769
rect 12139 34563 12173 34579
rect 11993 34529 12139 34563
rect 12139 34513 12173 34529
rect 55077 34563 55111 34579
rect 55111 34529 55257 34563
rect 55077 34513 55111 34529
rect 12139 34013 12173 34029
rect 11993 33979 12139 34013
rect 12139 33963 12173 33979
rect 55077 34013 55111 34029
rect 55111 33979 55257 34013
rect 55077 33963 55111 33979
rect 12139 33773 12173 33789
rect 11993 33739 12139 33773
rect 12139 33723 12173 33739
rect 55077 33773 55111 33789
rect 55111 33739 55257 33773
rect 55077 33723 55111 33739
rect 12139 33223 12173 33239
rect 11993 33189 12139 33223
rect 12139 33173 12173 33189
rect 55077 33223 55111 33239
rect 55111 33189 55257 33223
rect 55077 33173 55111 33189
rect 12139 32983 12173 32999
rect 11993 32949 12139 32983
rect 12139 32933 12173 32949
rect 55077 32983 55111 32999
rect 55111 32949 55257 32983
rect 55077 32933 55111 32949
rect 12139 32433 12173 32449
rect 11993 32399 12139 32433
rect 12139 32383 12173 32399
rect 55077 32433 55111 32449
rect 55111 32399 55257 32433
rect 55077 32383 55111 32399
rect 12139 32193 12173 32209
rect 11993 32159 12139 32193
rect 12139 32143 12173 32159
rect 55077 32193 55111 32209
rect 55111 32159 55257 32193
rect 55077 32143 55111 32159
rect 12139 31643 12173 31659
rect 11993 31609 12139 31643
rect 12139 31593 12173 31609
rect 55077 31643 55111 31659
rect 55111 31609 55257 31643
rect 55077 31593 55111 31609
rect 12139 31403 12173 31419
rect 11993 31369 12139 31403
rect 12139 31353 12173 31369
rect 55077 31403 55111 31419
rect 55111 31369 55257 31403
rect 55077 31353 55111 31369
rect 12139 30853 12173 30869
rect 11993 30819 12139 30853
rect 12139 30803 12173 30819
rect 55077 30853 55111 30869
rect 55111 30819 55257 30853
rect 55077 30803 55111 30819
rect 12139 30613 12173 30629
rect 11993 30579 12139 30613
rect 12139 30563 12173 30579
rect 55077 30613 55111 30629
rect 55111 30579 55257 30613
rect 55077 30563 55111 30579
rect 12139 30063 12173 30079
rect 11993 30029 12139 30063
rect 12139 30013 12173 30029
rect 55077 30063 55111 30079
rect 55111 30029 55257 30063
rect 55077 30013 55111 30029
rect 12139 29823 12173 29839
rect 11993 29789 12139 29823
rect 12139 29773 12173 29789
rect 55077 29823 55111 29839
rect 55111 29789 55257 29823
rect 55077 29773 55111 29789
rect 12139 29273 12173 29289
rect 11993 29239 12139 29273
rect 12139 29223 12173 29239
rect 55077 29273 55111 29289
rect 55111 29239 55257 29273
rect 55077 29223 55111 29239
rect 12139 29033 12173 29049
rect 11993 28999 12139 29033
rect 12139 28983 12173 28999
rect 55077 29033 55111 29049
rect 55111 28999 55257 29033
rect 55077 28983 55111 28999
rect 12139 28483 12173 28499
rect 11993 28449 12139 28483
rect 12139 28433 12173 28449
rect 55077 28483 55111 28499
rect 55111 28449 55257 28483
rect 55077 28433 55111 28449
rect 12139 28243 12173 28259
rect 11993 28209 12139 28243
rect 12139 28193 12173 28209
rect 55077 28243 55111 28259
rect 55111 28209 55257 28243
rect 55077 28193 55111 28209
rect 12139 27693 12173 27709
rect 11993 27659 12139 27693
rect 12139 27643 12173 27659
rect 55077 27693 55111 27709
rect 55111 27659 55257 27693
rect 55077 27643 55111 27659
rect 12139 27453 12173 27469
rect 11993 27419 12139 27453
rect 12139 27403 12173 27419
rect 55077 27453 55111 27469
rect 55111 27419 55257 27453
rect 55077 27403 55111 27419
rect 12139 26903 12173 26919
rect 11993 26869 12139 26903
rect 12139 26853 12173 26869
rect 55077 26903 55111 26919
rect 55111 26869 55257 26903
rect 55077 26853 55111 26869
rect 12139 26663 12173 26679
rect 11993 26629 12139 26663
rect 12139 26613 12173 26629
rect 55077 26663 55111 26679
rect 55111 26629 55257 26663
rect 55077 26613 55111 26629
rect 12139 26113 12173 26129
rect 11993 26079 12139 26113
rect 12139 26063 12173 26079
rect 55077 26113 55111 26129
rect 55111 26079 55257 26113
rect 55077 26063 55111 26079
rect 12139 25873 12173 25889
rect 11993 25839 12139 25873
rect 12139 25823 12173 25839
rect 55077 25873 55111 25889
rect 55111 25839 55257 25873
rect 55077 25823 55111 25839
rect 12139 25323 12173 25339
rect 11993 25289 12139 25323
rect 12139 25273 12173 25289
rect 55077 25323 55111 25339
rect 55111 25289 55257 25323
rect 55077 25273 55111 25289
rect 12139 25083 12173 25099
rect 11993 25049 12139 25083
rect 12139 25033 12173 25049
rect 55077 25083 55111 25099
rect 55111 25049 55257 25083
rect 55077 25033 55111 25049
rect 12139 24533 12173 24549
rect 11993 24499 12139 24533
rect 12139 24483 12173 24499
rect 55077 24533 55111 24549
rect 55111 24499 55257 24533
rect 55077 24483 55111 24499
rect 12139 24293 12173 24309
rect 11993 24259 12139 24293
rect 12139 24243 12173 24259
rect 55077 24293 55111 24309
rect 55111 24259 55257 24293
rect 55077 24243 55111 24259
rect 12139 23743 12173 23759
rect 11993 23709 12139 23743
rect 12139 23693 12173 23709
rect 55077 23743 55111 23759
rect 55111 23709 55257 23743
rect 55077 23693 55111 23709
rect 12139 23503 12173 23519
rect 11993 23469 12139 23503
rect 12139 23453 12173 23469
rect 55077 23503 55111 23519
rect 55111 23469 55257 23503
rect 55077 23453 55111 23469
rect 12139 22953 12173 22969
rect 11993 22919 12139 22953
rect 12139 22903 12173 22919
rect 55077 22953 55111 22969
rect 55111 22919 55257 22953
rect 55077 22903 55111 22919
rect 12139 22713 12173 22729
rect 11993 22679 12139 22713
rect 12139 22663 12173 22679
rect 55077 22713 55111 22729
rect 55111 22679 55257 22713
rect 55077 22663 55111 22679
rect 12139 22163 12173 22179
rect 11993 22129 12139 22163
rect 12139 22113 12173 22129
rect 55077 22163 55111 22179
rect 55111 22129 55257 22163
rect 55077 22113 55111 22129
rect 12139 21923 12173 21939
rect 11993 21889 12139 21923
rect 12139 21873 12173 21889
rect 55077 21923 55111 21939
rect 55111 21889 55257 21923
rect 55077 21873 55111 21889
rect 12139 21373 12173 21389
rect 11993 21339 12139 21373
rect 12139 21323 12173 21339
rect 55077 21373 55111 21389
rect 55111 21339 55257 21373
rect 55077 21323 55111 21339
rect 12139 21133 12173 21149
rect 11993 21099 12139 21133
rect 12139 21083 12173 21099
rect 55077 21133 55111 21149
rect 55111 21099 55257 21133
rect 55077 21083 55111 21099
rect 12139 20583 12173 20599
rect 11993 20549 12139 20583
rect 12139 20533 12173 20549
rect 55077 20583 55111 20599
rect 55111 20549 55257 20583
rect 55077 20533 55111 20549
rect 12139 20343 12173 20359
rect 11993 20309 12139 20343
rect 12139 20293 12173 20309
rect 55077 20343 55111 20359
rect 55111 20309 55257 20343
rect 55077 20293 55111 20309
rect 12139 19793 12173 19809
rect 11993 19759 12139 19793
rect 12139 19743 12173 19759
rect 55077 19793 55111 19809
rect 55111 19759 55257 19793
rect 55077 19743 55111 19759
rect 12139 19553 12173 19569
rect 11993 19519 12139 19553
rect 12139 19503 12173 19519
rect 55077 19553 55111 19569
rect 55111 19519 55257 19553
rect 55077 19503 55111 19519
rect 12139 19003 12173 19019
rect 11993 18969 12139 19003
rect 12139 18953 12173 18969
rect 55077 19003 55111 19019
rect 55111 18969 55257 19003
rect 55077 18953 55111 18969
rect 12139 18763 12173 18779
rect 11993 18729 12139 18763
rect 12139 18713 12173 18729
rect 55077 18763 55111 18779
rect 55111 18729 55257 18763
rect 55077 18713 55111 18729
rect 12139 18213 12173 18229
rect 11993 18179 12139 18213
rect 12139 18163 12173 18179
rect 55077 18213 55111 18229
rect 55111 18179 55257 18213
rect 55077 18163 55111 18179
rect 12139 17973 12173 17989
rect 11993 17939 12139 17973
rect 12139 17923 12173 17939
rect 55077 17973 55111 17989
rect 55111 17939 55257 17973
rect 55077 17923 55111 17939
rect 12139 17423 12173 17439
rect 11993 17389 12139 17423
rect 12139 17373 12173 17389
rect 55077 17423 55111 17439
rect 55111 17389 55257 17423
rect 55077 17373 55111 17389
rect 12139 17183 12173 17199
rect 11993 17149 12139 17183
rect 12139 17133 12173 17149
rect 55077 17183 55111 17199
rect 55111 17149 55257 17183
rect 55077 17133 55111 17149
rect 12139 16633 12173 16649
rect 11993 16599 12139 16633
rect 12139 16583 12173 16599
rect 55077 16633 55111 16649
rect 55111 16599 55257 16633
rect 55077 16583 55111 16599
rect 12139 16393 12173 16409
rect 11993 16359 12139 16393
rect 12139 16343 12173 16359
rect 55077 16393 55111 16409
rect 55111 16359 55257 16393
rect 55077 16343 55111 16359
rect 12139 15843 12173 15859
rect 11993 15809 12139 15843
rect 12139 15793 12173 15809
rect 55077 15843 55111 15859
rect 55111 15809 55257 15843
rect 55077 15793 55111 15809
rect 12139 15603 12173 15619
rect 11993 15569 12139 15603
rect 12139 15553 12173 15569
rect 55077 15603 55111 15619
rect 55111 15569 55257 15603
rect 55077 15553 55111 15569
rect 12139 15053 12173 15069
rect 11993 15019 12139 15053
rect 12139 15003 12173 15019
rect 55077 15053 55111 15069
rect 55111 15019 55257 15053
rect 55077 15003 55111 15019
rect 12139 14813 12173 14829
rect 11993 14779 12139 14813
rect 12139 14763 12173 14779
rect 55077 14813 55111 14829
rect 55111 14779 55257 14813
rect 55077 14763 55111 14779
rect 12139 14263 12173 14279
rect 11993 14229 12139 14263
rect 12139 14213 12173 14229
rect 55077 14263 55111 14279
rect 55111 14229 55257 14263
rect 55077 14213 55111 14229
rect 12139 14023 12173 14039
rect 11993 13989 12139 14023
rect 12139 13973 12173 13989
rect 55077 14023 55111 14039
rect 55111 13989 55257 14023
rect 55077 13973 55111 13989
rect 12139 13473 12173 13489
rect 11993 13439 12139 13473
rect 12139 13423 12173 13439
rect 55077 13473 55111 13489
rect 55111 13439 55257 13473
rect 55077 13423 55111 13439
rect 12139 13233 12173 13249
rect 11993 13199 12139 13233
rect 12139 13183 12173 13199
rect 55077 13233 55111 13249
rect 55111 13199 55257 13233
rect 55077 13183 55111 13199
rect 12139 12683 12173 12699
rect 11993 12649 12139 12683
rect 12139 12633 12173 12649
rect 55077 12683 55111 12699
rect 55111 12649 55257 12683
rect 55077 12633 55111 12649
rect 12139 12443 12173 12459
rect 11993 12409 12139 12443
rect 12139 12393 12173 12409
rect 55077 12443 55111 12459
rect 55111 12409 55257 12443
rect 55077 12393 55111 12409
rect 12139 11893 12173 11909
rect 11993 11859 12139 11893
rect 12139 11843 12173 11859
rect 55077 11893 55111 11909
rect 55111 11859 55257 11893
rect 55077 11843 55111 11859
rect 12139 11653 12173 11669
rect 11993 11619 12139 11653
rect 12139 11603 12173 11619
rect 55077 11653 55111 11669
rect 55111 11619 55257 11653
rect 55077 11603 55111 11619
rect 12139 11103 12173 11119
rect 11993 11069 12139 11103
rect 12139 11053 12173 11069
rect 55077 11103 55111 11119
rect 55111 11069 55257 11103
rect 55077 11053 55111 11069
rect 12139 10863 12173 10879
rect 11993 10829 12139 10863
rect 12139 10813 12173 10829
rect 55077 10863 55111 10879
rect 55111 10829 55257 10863
rect 55077 10813 55111 10829
rect 12139 10313 12173 10329
rect 11993 10279 12139 10313
rect 12139 10263 12173 10279
rect 55077 10313 55111 10329
rect 55111 10279 55257 10313
rect 55077 10263 55111 10279
rect 12139 10073 12173 10089
rect 11993 10039 12139 10073
rect 12139 10023 12173 10039
rect 6740 7652 6774 7668
rect 6740 7602 6774 7618
rect 7139 6945 7173 6961
rect 7139 6895 7173 6911
rect 6740 6238 6774 6254
rect 6740 6188 6774 6204
rect 7139 5531 7173 5547
rect 6053 5459 6087 5493
rect 7139 5481 7173 5497
rect 6740 4824 6774 4840
rect 6740 4774 6774 4790
<< viali >>
rect 60352 66088 60386 66122
rect 59953 65381 59987 65415
rect 60352 64674 60386 64708
rect 59953 63967 59987 64001
rect 60352 63260 60386 63294
rect 55077 60839 55111 60873
rect 12139 60599 12173 60633
rect 55077 60599 55111 60633
rect 12139 60049 12173 60083
rect 55077 60049 55111 60083
rect 12139 59809 12173 59843
rect 55077 59809 55111 59843
rect 12139 59259 12173 59293
rect 55077 59259 55111 59293
rect 12139 59019 12173 59053
rect 55077 59019 55111 59053
rect 12139 58469 12173 58503
rect 55077 58469 55111 58503
rect 12139 58229 12173 58263
rect 55077 58229 55111 58263
rect 12139 57679 12173 57713
rect 55077 57679 55111 57713
rect 12139 57439 12173 57473
rect 55077 57439 55111 57473
rect 12139 56889 12173 56923
rect 55077 56889 55111 56923
rect 12139 56649 12173 56683
rect 55077 56649 55111 56683
rect 12139 56099 12173 56133
rect 55077 56099 55111 56133
rect 12139 55859 12173 55893
rect 55077 55859 55111 55893
rect 12139 55309 12173 55343
rect 55077 55309 55111 55343
rect 12139 55069 12173 55103
rect 55077 55069 55111 55103
rect 12139 54519 12173 54553
rect 55077 54519 55111 54553
rect 12139 54279 12173 54313
rect 55077 54279 55111 54313
rect 12139 53729 12173 53763
rect 55077 53729 55111 53763
rect 12139 53489 12173 53523
rect 55077 53489 55111 53523
rect 12139 52939 12173 52973
rect 55077 52939 55111 52973
rect 12139 52699 12173 52733
rect 55077 52699 55111 52733
rect 12139 52149 12173 52183
rect 55077 52149 55111 52183
rect 12139 51909 12173 51943
rect 55077 51909 55111 51943
rect 12139 51359 12173 51393
rect 55077 51359 55111 51393
rect 12139 51119 12173 51153
rect 55077 51119 55111 51153
rect 12139 50569 12173 50603
rect 55077 50569 55111 50603
rect 12139 50329 12173 50363
rect 55077 50329 55111 50363
rect 12139 49779 12173 49813
rect 55077 49779 55111 49813
rect 12139 49539 12173 49573
rect 55077 49539 55111 49573
rect 12139 48989 12173 49023
rect 55077 48989 55111 49023
rect 12139 48749 12173 48783
rect 55077 48749 55111 48783
rect 12139 48199 12173 48233
rect 55077 48199 55111 48233
rect 12139 47959 12173 47993
rect 55077 47959 55111 47993
rect 12139 47409 12173 47443
rect 55077 47409 55111 47443
rect 12139 47169 12173 47203
rect 55077 47169 55111 47203
rect 12139 46619 12173 46653
rect 55077 46619 55111 46653
rect 12139 46379 12173 46413
rect 55077 46379 55111 46413
rect 12139 45829 12173 45863
rect 55077 45829 55111 45863
rect 12139 45589 12173 45623
rect 55077 45589 55111 45623
rect 12139 45039 12173 45073
rect 55077 45039 55111 45073
rect 12139 44799 12173 44833
rect 55077 44799 55111 44833
rect 12139 44249 12173 44283
rect 55077 44249 55111 44283
rect 12139 44009 12173 44043
rect 55077 44009 55111 44043
rect 12139 43459 12173 43493
rect 55077 43459 55111 43493
rect 12139 43219 12173 43253
rect 55077 43219 55111 43253
rect 12139 42669 12173 42703
rect 55077 42669 55111 42703
rect 12139 42429 12173 42463
rect 55077 42429 55111 42463
rect 12139 41879 12173 41913
rect 55077 41879 55111 41913
rect 12139 41639 12173 41673
rect 55077 41639 55111 41673
rect 12139 41089 12173 41123
rect 55077 41089 55111 41123
rect 12139 40849 12173 40883
rect 55077 40849 55111 40883
rect 12139 40299 12173 40333
rect 55077 40299 55111 40333
rect 12139 40059 12173 40093
rect 55077 40059 55111 40093
rect 12139 39509 12173 39543
rect 55077 39509 55111 39543
rect 12139 39269 12173 39303
rect 55077 39269 55111 39303
rect 12139 38719 12173 38753
rect 55077 38719 55111 38753
rect 12139 38479 12173 38513
rect 55077 38479 55111 38513
rect 12139 37929 12173 37963
rect 55077 37929 55111 37963
rect 12139 37689 12173 37723
rect 55077 37689 55111 37723
rect 12139 37139 12173 37173
rect 55077 37139 55111 37173
rect 12139 36899 12173 36933
rect 55077 36899 55111 36933
rect 12139 36349 12173 36383
rect 55077 36349 55111 36383
rect 12139 36109 12173 36143
rect 55077 36109 55111 36143
rect 12139 35559 12173 35593
rect 55077 35559 55111 35593
rect 12139 35319 12173 35353
rect 55077 35319 55111 35353
rect 12139 34769 12173 34803
rect 55077 34769 55111 34803
rect 12139 34529 12173 34563
rect 55077 34529 55111 34563
rect 12139 33979 12173 34013
rect 55077 33979 55111 34013
rect 12139 33739 12173 33773
rect 55077 33739 55111 33773
rect 12139 33189 12173 33223
rect 55077 33189 55111 33223
rect 12139 32949 12173 32983
rect 55077 32949 55111 32983
rect 12139 32399 12173 32433
rect 55077 32399 55111 32433
rect 12139 32159 12173 32193
rect 55077 32159 55111 32193
rect 12139 31609 12173 31643
rect 55077 31609 55111 31643
rect 12139 31369 12173 31403
rect 55077 31369 55111 31403
rect 12139 30819 12173 30853
rect 55077 30819 55111 30853
rect 12139 30579 12173 30613
rect 55077 30579 55111 30613
rect 12139 30029 12173 30063
rect 55077 30029 55111 30063
rect 12139 29789 12173 29823
rect 55077 29789 55111 29823
rect 12139 29239 12173 29273
rect 55077 29239 55111 29273
rect 12139 28999 12173 29033
rect 55077 28999 55111 29033
rect 12139 28449 12173 28483
rect 55077 28449 55111 28483
rect 12139 28209 12173 28243
rect 55077 28209 55111 28243
rect 12139 27659 12173 27693
rect 55077 27659 55111 27693
rect 12139 27419 12173 27453
rect 55077 27419 55111 27453
rect 12139 26869 12173 26903
rect 55077 26869 55111 26903
rect 12139 26629 12173 26663
rect 55077 26629 55111 26663
rect 12139 26079 12173 26113
rect 55077 26079 55111 26113
rect 12139 25839 12173 25873
rect 55077 25839 55111 25873
rect 12139 25289 12173 25323
rect 55077 25289 55111 25323
rect 12139 25049 12173 25083
rect 55077 25049 55111 25083
rect 12139 24499 12173 24533
rect 55077 24499 55111 24533
rect 12139 24259 12173 24293
rect 55077 24259 55111 24293
rect 12139 23709 12173 23743
rect 55077 23709 55111 23743
rect 12139 23469 12173 23503
rect 55077 23469 55111 23503
rect 12139 22919 12173 22953
rect 55077 22919 55111 22953
rect 12139 22679 12173 22713
rect 55077 22679 55111 22713
rect 12139 22129 12173 22163
rect 55077 22129 55111 22163
rect 12139 21889 12173 21923
rect 55077 21889 55111 21923
rect 12139 21339 12173 21373
rect 55077 21339 55111 21373
rect 12139 21099 12173 21133
rect 55077 21099 55111 21133
rect 12139 20549 12173 20583
rect 55077 20549 55111 20583
rect 12139 20309 12173 20343
rect 55077 20309 55111 20343
rect 12139 19759 12173 19793
rect 55077 19759 55111 19793
rect 12139 19519 12173 19553
rect 55077 19519 55111 19553
rect 12139 18969 12173 19003
rect 55077 18969 55111 19003
rect 12139 18729 12173 18763
rect 55077 18729 55111 18763
rect 12139 18179 12173 18213
rect 55077 18179 55111 18213
rect 12139 17939 12173 17973
rect 55077 17939 55111 17973
rect 12139 17389 12173 17423
rect 55077 17389 55111 17423
rect 12139 17149 12173 17183
rect 55077 17149 55111 17183
rect 12139 16599 12173 16633
rect 55077 16599 55111 16633
rect 12139 16359 12173 16393
rect 55077 16359 55111 16393
rect 12139 15809 12173 15843
rect 55077 15809 55111 15843
rect 12139 15569 12173 15603
rect 55077 15569 55111 15603
rect 12139 15019 12173 15053
rect 55077 15019 55111 15053
rect 12139 14779 12173 14813
rect 55077 14779 55111 14813
rect 12139 14229 12173 14263
rect 55077 14229 55111 14263
rect 12139 13989 12173 14023
rect 55077 13989 55111 14023
rect 12139 13439 12173 13473
rect 55077 13439 55111 13473
rect 12139 13199 12173 13233
rect 55077 13199 55111 13233
rect 12139 12649 12173 12683
rect 55077 12649 55111 12683
rect 12139 12409 12173 12443
rect 55077 12409 55111 12443
rect 12139 11859 12173 11893
rect 55077 11859 55111 11893
rect 12139 11619 12173 11653
rect 55077 11619 55111 11653
rect 12139 11069 12173 11103
rect 55077 11069 55111 11103
rect 12139 10829 12173 10863
rect 55077 10829 55111 10863
rect 12139 10279 12173 10313
rect 55077 10279 55111 10313
rect 12139 10039 12173 10073
rect 6740 7618 6774 7652
rect 7139 6911 7173 6945
rect 6740 6204 6774 6238
rect 7139 5497 7173 5531
rect 6740 4790 6774 4824
<< metal1 >>
rect 13761 66974 13807 67228
rect 15009 66974 15055 67228
rect 16257 66974 16303 67228
rect 17505 66974 17551 67228
rect 18753 66974 18799 67228
rect 20001 66974 20047 67228
rect 21249 66974 21295 67228
rect 22497 66974 22543 67228
rect 23745 66974 23791 67228
rect 24993 66974 25039 67228
rect 26241 66974 26287 67228
rect 27489 66974 27535 67228
rect 28737 66974 28783 67228
rect 29985 66974 30031 67228
rect 31233 66974 31279 67228
rect 32481 66974 32527 67228
rect 33729 66974 33775 67228
rect 34977 66974 35023 67228
rect 36225 66974 36271 67228
rect 37473 66974 37519 67228
rect 38721 66974 38767 67228
rect 39969 66974 40015 67228
rect 41217 66974 41263 67228
rect 42465 66974 42511 67228
rect 43713 66974 43759 67228
rect 44961 66974 45007 67228
rect 46209 66974 46255 67228
rect 47457 66974 47503 67228
rect 48705 66974 48751 67228
rect 49953 66974 49999 67228
rect 51201 66974 51247 67228
rect 52449 66974 52495 67228
rect 60337 66079 60343 66131
rect 60395 66079 60401 66131
rect 59938 65372 59944 65424
rect 59996 65372 60002 65424
rect 60337 64665 60343 64717
rect 60395 64665 60401 64717
rect 59938 63958 59944 64010
rect 59996 63958 60002 64010
rect 60337 63251 60343 63303
rect 60395 63251 60401 63303
rect 53641 62630 53647 62682
rect 53699 62630 53705 62682
rect 53659 62532 53687 62630
rect 13723 61666 13751 61778
rect 14187 61666 14215 61778
rect 13723 61638 13983 61666
rect 13955 61526 13983 61638
rect 14027 61638 14215 61666
rect 14347 61666 14375 61778
rect 14811 61666 14839 61778
rect 14347 61638 14535 61666
rect 14027 61526 14055 61638
rect 14507 61526 14535 61638
rect 14579 61638 14839 61666
rect 14971 61666 14999 61778
rect 15435 61666 15463 61778
rect 14971 61638 15231 61666
rect 14579 61526 14607 61638
rect 15203 61526 15231 61638
rect 15275 61638 15463 61666
rect 15595 61666 15623 61778
rect 16059 61666 16087 61778
rect 15595 61638 15783 61666
rect 15275 61526 15303 61638
rect 15755 61526 15783 61638
rect 15827 61638 16087 61666
rect 16219 61666 16247 61778
rect 16683 61666 16711 61778
rect 16219 61638 16479 61666
rect 15827 61526 15855 61638
rect 16451 61526 16479 61638
rect 16523 61638 16711 61666
rect 16843 61666 16871 61778
rect 17307 61666 17335 61778
rect 16843 61638 17031 61666
rect 16523 61526 16551 61638
rect 17003 61526 17031 61638
rect 17075 61638 17335 61666
rect 17467 61666 17495 61778
rect 17931 61666 17959 61778
rect 17467 61638 17727 61666
rect 17075 61526 17103 61638
rect 17699 61526 17727 61638
rect 17771 61638 17959 61666
rect 18091 61666 18119 61778
rect 18555 61666 18583 61778
rect 18091 61638 18279 61666
rect 17771 61526 17799 61638
rect 18251 61526 18279 61638
rect 18323 61638 18583 61666
rect 18715 61666 18743 61778
rect 19179 61666 19207 61778
rect 18715 61638 18975 61666
rect 18323 61526 18351 61638
rect 18947 61526 18975 61638
rect 19019 61638 19207 61666
rect 19339 61666 19367 61778
rect 19803 61666 19831 61778
rect 19339 61638 19527 61666
rect 19019 61526 19047 61638
rect 19499 61526 19527 61638
rect 19571 61638 19831 61666
rect 19963 61666 19991 61778
rect 20427 61666 20455 61778
rect 19963 61638 20223 61666
rect 19571 61526 19599 61638
rect 20195 61526 20223 61638
rect 20267 61638 20455 61666
rect 20587 61666 20615 61778
rect 21051 61666 21079 61778
rect 20587 61638 20775 61666
rect 20267 61526 20295 61638
rect 20747 61526 20775 61638
rect 20819 61638 21079 61666
rect 21211 61666 21239 61778
rect 21675 61666 21703 61778
rect 21211 61638 21471 61666
rect 20819 61526 20847 61638
rect 21443 61526 21471 61638
rect 21515 61638 21703 61666
rect 21835 61666 21863 61778
rect 22299 61666 22327 61778
rect 21835 61638 22023 61666
rect 21515 61526 21543 61638
rect 21995 61526 22023 61638
rect 22067 61638 22327 61666
rect 22459 61666 22487 61778
rect 22923 61666 22951 61778
rect 22459 61638 22719 61666
rect 22067 61526 22095 61638
rect 22691 61526 22719 61638
rect 22763 61638 22951 61666
rect 23083 61666 23111 61778
rect 23547 61666 23575 61778
rect 23083 61638 23271 61666
rect 22763 61526 22791 61638
rect 23243 61526 23271 61638
rect 23315 61638 23575 61666
rect 23707 61666 23735 61778
rect 24171 61666 24199 61778
rect 23707 61638 23967 61666
rect 23315 61526 23343 61638
rect 23939 61526 23967 61638
rect 24011 61638 24199 61666
rect 24331 61666 24359 61778
rect 24795 61666 24823 61778
rect 24331 61638 24519 61666
rect 24011 61526 24039 61638
rect 24491 61526 24519 61638
rect 24563 61638 24823 61666
rect 24955 61666 24983 61778
rect 25419 61666 25447 61778
rect 24955 61638 25215 61666
rect 24563 61526 24591 61638
rect 25187 61526 25215 61638
rect 25259 61638 25447 61666
rect 25579 61666 25607 61778
rect 26043 61666 26071 61778
rect 25579 61638 25767 61666
rect 25259 61526 25287 61638
rect 25739 61526 25767 61638
rect 25811 61638 26071 61666
rect 26203 61666 26231 61778
rect 26667 61666 26695 61778
rect 26203 61638 26463 61666
rect 25811 61526 25839 61638
rect 26435 61526 26463 61638
rect 26507 61638 26695 61666
rect 26827 61666 26855 61778
rect 27291 61666 27319 61778
rect 26827 61638 27015 61666
rect 26507 61526 26535 61638
rect 26987 61526 27015 61638
rect 27059 61638 27319 61666
rect 27451 61666 27479 61778
rect 27915 61666 27943 61778
rect 27451 61638 27711 61666
rect 27059 61526 27087 61638
rect 27683 61526 27711 61638
rect 27755 61638 27943 61666
rect 28075 61666 28103 61778
rect 28539 61666 28567 61778
rect 28075 61638 28263 61666
rect 27755 61526 27783 61638
rect 28235 61526 28263 61638
rect 28307 61638 28567 61666
rect 28699 61666 28727 61778
rect 29163 61666 29191 61778
rect 28699 61638 28959 61666
rect 28307 61526 28335 61638
rect 28931 61526 28959 61638
rect 29003 61638 29191 61666
rect 29323 61666 29351 61778
rect 29787 61666 29815 61778
rect 29323 61638 29511 61666
rect 29003 61526 29031 61638
rect 29483 61526 29511 61638
rect 29555 61638 29815 61666
rect 29947 61666 29975 61778
rect 30411 61666 30439 61778
rect 29947 61638 30207 61666
rect 29555 61526 29583 61638
rect 30179 61526 30207 61638
rect 30251 61638 30439 61666
rect 30571 61666 30599 61778
rect 31035 61666 31063 61778
rect 30571 61638 30759 61666
rect 30251 61526 30279 61638
rect 30731 61526 30759 61638
rect 30803 61638 31063 61666
rect 31195 61666 31223 61778
rect 31659 61666 31687 61778
rect 31195 61638 31455 61666
rect 30803 61526 30831 61638
rect 31427 61526 31455 61638
rect 31499 61638 31687 61666
rect 31819 61666 31847 61778
rect 32283 61666 32311 61778
rect 31819 61638 32007 61666
rect 31499 61526 31527 61638
rect 31979 61526 32007 61638
rect 32051 61638 32311 61666
rect 32443 61666 32471 61778
rect 32907 61666 32935 61778
rect 32443 61638 32703 61666
rect 32051 61526 32079 61638
rect 32675 61526 32703 61638
rect 32747 61638 32935 61666
rect 33067 61666 33095 61778
rect 33531 61666 33559 61778
rect 33067 61638 33255 61666
rect 32747 61526 32775 61638
rect 33227 61526 33255 61638
rect 33299 61638 33559 61666
rect 33691 61666 33719 61778
rect 34155 61666 34183 61778
rect 33691 61638 33951 61666
rect 33299 61526 33327 61638
rect 33923 61526 33951 61638
rect 33995 61638 34183 61666
rect 34315 61666 34343 61778
rect 34779 61666 34807 61778
rect 34315 61638 34503 61666
rect 33995 61526 34023 61638
rect 34475 61526 34503 61638
rect 34547 61638 34807 61666
rect 34939 61666 34967 61778
rect 35403 61666 35431 61778
rect 34939 61638 35199 61666
rect 34547 61526 34575 61638
rect 35171 61526 35199 61638
rect 35243 61638 35431 61666
rect 35563 61666 35591 61778
rect 36027 61666 36055 61778
rect 35563 61638 35751 61666
rect 35243 61526 35271 61638
rect 35723 61526 35751 61638
rect 35795 61638 36055 61666
rect 36187 61666 36215 61778
rect 36651 61666 36679 61778
rect 36187 61638 36447 61666
rect 35795 61526 35823 61638
rect 36419 61526 36447 61638
rect 36491 61638 36679 61666
rect 36811 61666 36839 61778
rect 37275 61666 37303 61778
rect 36811 61638 36999 61666
rect 36491 61526 36519 61638
rect 36971 61526 36999 61638
rect 37043 61638 37303 61666
rect 37435 61666 37463 61778
rect 37899 61666 37927 61778
rect 37435 61638 37695 61666
rect 37043 61526 37071 61638
rect 37667 61526 37695 61638
rect 37739 61638 37927 61666
rect 38059 61666 38087 61778
rect 38523 61666 38551 61778
rect 38059 61638 38247 61666
rect 37739 61526 37767 61638
rect 38219 61526 38247 61638
rect 38291 61638 38551 61666
rect 38683 61666 38711 61778
rect 39147 61666 39175 61778
rect 38683 61638 38943 61666
rect 38291 61526 38319 61638
rect 38915 61526 38943 61638
rect 38987 61638 39175 61666
rect 39307 61666 39335 61778
rect 39771 61666 39799 61778
rect 39307 61638 39495 61666
rect 38987 61526 39015 61638
rect 39467 61526 39495 61638
rect 39539 61638 39799 61666
rect 39931 61666 39959 61778
rect 40395 61666 40423 61778
rect 39931 61638 40191 61666
rect 39539 61526 39567 61638
rect 40163 61526 40191 61638
rect 40235 61638 40423 61666
rect 40555 61666 40583 61778
rect 41019 61666 41047 61778
rect 40555 61638 40743 61666
rect 40235 61526 40263 61638
rect 40715 61526 40743 61638
rect 40787 61638 41047 61666
rect 41179 61666 41207 61778
rect 41643 61666 41671 61778
rect 41179 61638 41439 61666
rect 40787 61526 40815 61638
rect 41411 61526 41439 61638
rect 41483 61638 41671 61666
rect 41803 61666 41831 61778
rect 42267 61666 42295 61778
rect 41803 61638 41991 61666
rect 41483 61526 41511 61638
rect 41963 61526 41991 61638
rect 42035 61638 42295 61666
rect 42427 61666 42455 61778
rect 42891 61666 42919 61778
rect 42427 61638 42687 61666
rect 42035 61526 42063 61638
rect 42659 61526 42687 61638
rect 42731 61638 42919 61666
rect 43051 61666 43079 61778
rect 43515 61666 43543 61778
rect 43051 61638 43239 61666
rect 42731 61526 42759 61638
rect 43211 61526 43239 61638
rect 43283 61638 43543 61666
rect 43675 61666 43703 61778
rect 44139 61666 44167 61778
rect 43675 61638 43935 61666
rect 43283 61526 43311 61638
rect 43907 61526 43935 61638
rect 43979 61638 44167 61666
rect 44299 61666 44327 61778
rect 44763 61666 44791 61778
rect 44299 61638 44487 61666
rect 43979 61526 44007 61638
rect 44459 61526 44487 61638
rect 44531 61638 44791 61666
rect 44923 61666 44951 61778
rect 45387 61666 45415 61778
rect 44923 61638 45183 61666
rect 44531 61526 44559 61638
rect 45155 61526 45183 61638
rect 45227 61638 45415 61666
rect 45547 61666 45575 61778
rect 46011 61666 46039 61778
rect 45547 61638 45735 61666
rect 45227 61526 45255 61638
rect 45707 61526 45735 61638
rect 45779 61638 46039 61666
rect 46171 61666 46199 61778
rect 46635 61666 46663 61778
rect 46171 61638 46431 61666
rect 45779 61526 45807 61638
rect 46403 61526 46431 61638
rect 46475 61638 46663 61666
rect 46795 61666 46823 61778
rect 47259 61666 47287 61778
rect 46795 61638 46983 61666
rect 46475 61526 46503 61638
rect 46955 61526 46983 61638
rect 47027 61638 47287 61666
rect 47419 61666 47447 61778
rect 47883 61666 47911 61778
rect 47419 61638 47679 61666
rect 47027 61526 47055 61638
rect 47651 61526 47679 61638
rect 47723 61638 47911 61666
rect 48043 61666 48071 61778
rect 48507 61666 48535 61778
rect 48043 61638 48231 61666
rect 47723 61526 47751 61638
rect 48203 61526 48231 61638
rect 48275 61638 48535 61666
rect 48667 61666 48695 61778
rect 49131 61666 49159 61778
rect 48667 61638 48927 61666
rect 48275 61526 48303 61638
rect 48899 61526 48927 61638
rect 48971 61638 49159 61666
rect 49291 61666 49319 61778
rect 49755 61666 49783 61778
rect 49291 61638 49479 61666
rect 48971 61526 48999 61638
rect 49451 61526 49479 61638
rect 49523 61638 49783 61666
rect 49915 61666 49943 61778
rect 50379 61666 50407 61778
rect 49915 61638 50175 61666
rect 49523 61526 49551 61638
rect 50147 61526 50175 61638
rect 50219 61638 50407 61666
rect 50539 61666 50567 61778
rect 51003 61666 51031 61778
rect 50539 61638 50727 61666
rect 50219 61526 50247 61638
rect 50699 61526 50727 61638
rect 50771 61638 51031 61666
rect 51163 61666 51191 61778
rect 51627 61666 51655 61778
rect 51163 61638 51423 61666
rect 50771 61526 50799 61638
rect 51395 61526 51423 61638
rect 51467 61638 51655 61666
rect 51787 61666 51815 61778
rect 52251 61666 52279 61778
rect 51787 61638 51975 61666
rect 51467 61526 51495 61638
rect 51947 61526 51975 61638
rect 52019 61638 52279 61666
rect 52411 61666 52439 61778
rect 52875 61666 52903 61778
rect 52411 61638 52671 61666
rect 52019 61526 52047 61638
rect 52643 61526 52671 61638
rect 52715 61638 52903 61666
rect 53035 61666 53063 61778
rect 53499 61666 53527 61778
rect 53035 61638 53223 61666
rect 52715 61526 52743 61638
rect 53195 61526 53223 61638
rect 53267 61638 53527 61666
rect 53659 61666 53687 61778
rect 54123 61666 54151 61778
rect 53659 61638 53919 61666
rect 53267 61526 53295 61638
rect 53891 61526 53919 61638
rect 53963 61638 54151 61666
rect 53963 61526 53991 61638
rect 55062 60830 55068 60882
rect 55120 60830 55126 60882
rect 12124 60590 12130 60642
rect 12182 60590 12188 60642
rect 55062 60590 55068 60642
rect 55120 60590 55126 60642
rect 12124 60040 12130 60092
rect 12182 60040 12188 60092
rect 55062 60040 55068 60092
rect 55120 60040 55126 60092
rect 12124 59800 12130 59852
rect 12182 59800 12188 59852
rect 55062 59800 55068 59852
rect 55120 59800 55126 59852
rect 12124 59250 12130 59302
rect 12182 59250 12188 59302
rect 55062 59250 55068 59302
rect 55120 59250 55126 59302
rect 12124 59010 12130 59062
rect 12182 59010 12188 59062
rect 55062 59010 55068 59062
rect 55120 59010 55126 59062
rect 12124 58460 12130 58512
rect 12182 58460 12188 58512
rect 55062 58460 55068 58512
rect 55120 58460 55126 58512
rect 12124 58220 12130 58272
rect 12182 58220 12188 58272
rect 55062 58220 55068 58272
rect 55120 58220 55126 58272
rect 12124 57670 12130 57722
rect 12182 57670 12188 57722
rect 55062 57670 55068 57722
rect 55120 57670 55126 57722
rect 12124 57430 12130 57482
rect 12182 57430 12188 57482
rect 55062 57430 55068 57482
rect 55120 57430 55126 57482
rect 12124 56880 12130 56932
rect 12182 56880 12188 56932
rect 55062 56880 55068 56932
rect 55120 56880 55126 56932
rect 12124 56640 12130 56692
rect 12182 56640 12188 56692
rect 55062 56640 55068 56692
rect 55120 56640 55126 56692
rect 12124 56090 12130 56142
rect 12182 56090 12188 56142
rect 55062 56090 55068 56142
rect 55120 56090 55126 56142
rect 12124 55850 12130 55902
rect 12182 55850 12188 55902
rect 55062 55850 55068 55902
rect 55120 55850 55126 55902
rect 12124 55300 12130 55352
rect 12182 55300 12188 55352
rect 55062 55300 55068 55352
rect 55120 55300 55126 55352
rect 12124 55060 12130 55112
rect 12182 55060 12188 55112
rect 55062 55060 55068 55112
rect 55120 55060 55126 55112
rect 12124 54510 12130 54562
rect 12182 54510 12188 54562
rect 55062 54510 55068 54562
rect 55120 54510 55126 54562
rect 12124 54270 12130 54322
rect 12182 54270 12188 54322
rect 55062 54270 55068 54322
rect 55120 54270 55126 54322
rect 12124 53720 12130 53772
rect 12182 53720 12188 53772
rect 55062 53720 55068 53772
rect 55120 53720 55126 53772
rect 12124 53480 12130 53532
rect 12182 53480 12188 53532
rect 55062 53480 55068 53532
rect 55120 53480 55126 53532
rect 12124 52930 12130 52982
rect 12182 52930 12188 52982
rect 55062 52930 55068 52982
rect 55120 52930 55126 52982
rect 12124 52690 12130 52742
rect 12182 52690 12188 52742
rect 55062 52690 55068 52742
rect 55120 52690 55126 52742
rect 12124 52140 12130 52192
rect 12182 52140 12188 52192
rect 55062 52140 55068 52192
rect 55120 52140 55126 52192
rect 12124 51900 12130 51952
rect 12182 51900 12188 51952
rect 55062 51900 55068 51952
rect 55120 51900 55126 51952
rect 12124 51350 12130 51402
rect 12182 51350 12188 51402
rect 55062 51350 55068 51402
rect 55120 51350 55126 51402
rect 12124 51110 12130 51162
rect 12182 51110 12188 51162
rect 55062 51110 55068 51162
rect 55120 51110 55126 51162
rect 12124 50560 12130 50612
rect 12182 50560 12188 50612
rect 55062 50560 55068 50612
rect 55120 50560 55126 50612
rect 12124 50320 12130 50372
rect 12182 50320 12188 50372
rect 55062 50320 55068 50372
rect 55120 50320 55126 50372
rect 12124 49770 12130 49822
rect 12182 49770 12188 49822
rect 55062 49770 55068 49822
rect 55120 49770 55126 49822
rect 12124 49530 12130 49582
rect 12182 49530 12188 49582
rect 55062 49530 55068 49582
rect 55120 49530 55126 49582
rect 12124 48980 12130 49032
rect 12182 48980 12188 49032
rect 55062 48980 55068 49032
rect 55120 48980 55126 49032
rect 12124 48740 12130 48792
rect 12182 48740 12188 48792
rect 55062 48740 55068 48792
rect 55120 48740 55126 48792
rect 12124 48190 12130 48242
rect 12182 48190 12188 48242
rect 55062 48190 55068 48242
rect 55120 48190 55126 48242
rect 12124 47950 12130 48002
rect 12182 47950 12188 48002
rect 55062 47950 55068 48002
rect 55120 47950 55126 48002
rect 12124 47400 12130 47452
rect 12182 47400 12188 47452
rect 55062 47400 55068 47452
rect 55120 47400 55126 47452
rect 12124 47160 12130 47212
rect 12182 47160 12188 47212
rect 55062 47160 55068 47212
rect 55120 47160 55126 47212
rect 12124 46610 12130 46662
rect 12182 46610 12188 46662
rect 55062 46610 55068 46662
rect 55120 46610 55126 46662
rect 12124 46370 12130 46422
rect 12182 46370 12188 46422
rect 55062 46370 55068 46422
rect 55120 46370 55126 46422
rect 12124 45820 12130 45872
rect 12182 45820 12188 45872
rect 55062 45820 55068 45872
rect 55120 45820 55126 45872
rect 12124 45580 12130 45632
rect 12182 45580 12188 45632
rect 55062 45580 55068 45632
rect 55120 45580 55126 45632
rect 12124 45030 12130 45082
rect 12182 45030 12188 45082
rect 55062 45030 55068 45082
rect 55120 45030 55126 45082
rect 12124 44790 12130 44842
rect 12182 44790 12188 44842
rect 55062 44790 55068 44842
rect 55120 44790 55126 44842
rect 12124 44240 12130 44292
rect 12182 44240 12188 44292
rect 55062 44240 55068 44292
rect 55120 44240 55126 44292
rect 12124 44000 12130 44052
rect 12182 44000 12188 44052
rect 55062 44000 55068 44052
rect 55120 44000 55126 44052
rect 12124 43450 12130 43502
rect 12182 43450 12188 43502
rect 55062 43450 55068 43502
rect 55120 43450 55126 43502
rect 12124 43210 12130 43262
rect 12182 43210 12188 43262
rect 55062 43210 55068 43262
rect 55120 43210 55126 43262
rect 12124 42660 12130 42712
rect 12182 42660 12188 42712
rect 55062 42660 55068 42712
rect 55120 42660 55126 42712
rect 12124 42420 12130 42472
rect 12182 42420 12188 42472
rect 55062 42420 55068 42472
rect 55120 42420 55126 42472
rect 12124 41870 12130 41922
rect 12182 41870 12188 41922
rect 55062 41870 55068 41922
rect 55120 41870 55126 41922
rect 12124 41630 12130 41682
rect 12182 41630 12188 41682
rect 55062 41630 55068 41682
rect 55120 41630 55126 41682
rect 12124 41080 12130 41132
rect 12182 41080 12188 41132
rect 55062 41080 55068 41132
rect 55120 41080 55126 41132
rect 12124 40840 12130 40892
rect 12182 40840 12188 40892
rect 55062 40840 55068 40892
rect 55120 40840 55126 40892
rect 12124 40290 12130 40342
rect 12182 40290 12188 40342
rect 55062 40290 55068 40342
rect 55120 40290 55126 40342
rect 12124 40050 12130 40102
rect 12182 40050 12188 40102
rect 55062 40050 55068 40102
rect 55120 40050 55126 40102
rect 12124 39500 12130 39552
rect 12182 39500 12188 39552
rect 55062 39500 55068 39552
rect 55120 39500 55126 39552
rect 12124 39260 12130 39312
rect 12182 39260 12188 39312
rect 55062 39260 55068 39312
rect 55120 39260 55126 39312
rect 12124 38710 12130 38762
rect 12182 38710 12188 38762
rect 55062 38710 55068 38762
rect 55120 38710 55126 38762
rect 12124 38470 12130 38522
rect 12182 38470 12188 38522
rect 55062 38470 55068 38522
rect 55120 38470 55126 38522
rect 12124 37920 12130 37972
rect 12182 37920 12188 37972
rect 55062 37920 55068 37972
rect 55120 37920 55126 37972
rect 12124 37680 12130 37732
rect 12182 37680 12188 37732
rect 55062 37680 55068 37732
rect 55120 37680 55126 37732
rect 12124 37130 12130 37182
rect 12182 37130 12188 37182
rect 55062 37130 55068 37182
rect 55120 37130 55126 37182
rect 12124 36890 12130 36942
rect 12182 36890 12188 36942
rect 55062 36890 55068 36942
rect 55120 36890 55126 36942
rect 12124 36340 12130 36392
rect 12182 36340 12188 36392
rect 55062 36340 55068 36392
rect 55120 36340 55126 36392
rect 12124 36100 12130 36152
rect 12182 36100 12188 36152
rect 55062 36100 55068 36152
rect 55120 36100 55126 36152
rect 12124 35550 12130 35602
rect 12182 35550 12188 35602
rect 55062 35550 55068 35602
rect 55120 35550 55126 35602
rect 12124 35310 12130 35362
rect 12182 35310 12188 35362
rect 55062 35310 55068 35362
rect 55120 35310 55126 35362
rect 12124 34760 12130 34812
rect 12182 34760 12188 34812
rect 55062 34760 55068 34812
rect 55120 34760 55126 34812
rect 12124 34520 12130 34572
rect 12182 34520 12188 34572
rect 55062 34520 55068 34572
rect 55120 34520 55126 34572
rect 12124 33970 12130 34022
rect 12182 33970 12188 34022
rect 55062 33970 55068 34022
rect 55120 33970 55126 34022
rect 12124 33730 12130 33782
rect 12182 33730 12188 33782
rect 55062 33730 55068 33782
rect 55120 33730 55126 33782
rect 12124 33180 12130 33232
rect 12182 33180 12188 33232
rect 55062 33180 55068 33232
rect 55120 33180 55126 33232
rect 12124 32940 12130 32992
rect 12182 32940 12188 32992
rect 55062 32940 55068 32992
rect 55120 32940 55126 32992
rect 12124 32390 12130 32442
rect 12182 32390 12188 32442
rect 55062 32390 55068 32442
rect 55120 32390 55126 32442
rect 12124 32150 12130 32202
rect 12182 32150 12188 32202
rect 55062 32150 55068 32202
rect 55120 32150 55126 32202
rect 12124 31600 12130 31652
rect 12182 31600 12188 31652
rect 55062 31600 55068 31652
rect 55120 31600 55126 31652
rect 12124 31360 12130 31412
rect 12182 31360 12188 31412
rect 55062 31360 55068 31412
rect 55120 31360 55126 31412
rect 12124 30810 12130 30862
rect 12182 30810 12188 30862
rect 55062 30810 55068 30862
rect 55120 30810 55126 30862
rect 12124 30570 12130 30622
rect 12182 30570 12188 30622
rect 55062 30570 55068 30622
rect 55120 30570 55126 30622
rect 12124 30020 12130 30072
rect 12182 30020 12188 30072
rect 55062 30020 55068 30072
rect 55120 30020 55126 30072
rect 12124 29780 12130 29832
rect 12182 29780 12188 29832
rect 55062 29780 55068 29832
rect 55120 29780 55126 29832
rect 12124 29230 12130 29282
rect 12182 29230 12188 29282
rect 55062 29230 55068 29282
rect 55120 29230 55126 29282
rect 12124 28990 12130 29042
rect 12182 28990 12188 29042
rect 55062 28990 55068 29042
rect 55120 28990 55126 29042
rect 12124 28440 12130 28492
rect 12182 28440 12188 28492
rect 55062 28440 55068 28492
rect 55120 28440 55126 28492
rect 12124 28200 12130 28252
rect 12182 28200 12188 28252
rect 55062 28200 55068 28252
rect 55120 28200 55126 28252
rect 12124 27650 12130 27702
rect 12182 27650 12188 27702
rect 55062 27650 55068 27702
rect 55120 27650 55126 27702
rect 12124 27410 12130 27462
rect 12182 27410 12188 27462
rect 55062 27410 55068 27462
rect 55120 27410 55126 27462
rect 12124 26860 12130 26912
rect 12182 26860 12188 26912
rect 55062 26860 55068 26912
rect 55120 26860 55126 26912
rect 12124 26620 12130 26672
rect 12182 26620 12188 26672
rect 55062 26620 55068 26672
rect 55120 26620 55126 26672
rect 12124 26070 12130 26122
rect 12182 26070 12188 26122
rect 55062 26070 55068 26122
rect 55120 26070 55126 26122
rect 12124 25830 12130 25882
rect 12182 25830 12188 25882
rect 55062 25830 55068 25882
rect 55120 25830 55126 25882
rect 12124 25280 12130 25332
rect 12182 25280 12188 25332
rect 55062 25280 55068 25332
rect 55120 25280 55126 25332
rect 12124 25040 12130 25092
rect 12182 25040 12188 25092
rect 55062 25040 55068 25092
rect 55120 25040 55126 25092
rect 12124 24490 12130 24542
rect 12182 24490 12188 24542
rect 55062 24490 55068 24542
rect 55120 24490 55126 24542
rect 12124 24250 12130 24302
rect 12182 24250 12188 24302
rect 55062 24250 55068 24302
rect 55120 24250 55126 24302
rect 12124 23700 12130 23752
rect 12182 23700 12188 23752
rect 55062 23700 55068 23752
rect 55120 23700 55126 23752
rect 12124 23460 12130 23512
rect 12182 23460 12188 23512
rect 55062 23460 55068 23512
rect 55120 23460 55126 23512
rect 12124 22910 12130 22962
rect 12182 22910 12188 22962
rect 55062 22910 55068 22962
rect 55120 22910 55126 22962
rect 12124 22670 12130 22722
rect 12182 22670 12188 22722
rect 55062 22670 55068 22722
rect 55120 22670 55126 22722
rect 12124 22120 12130 22172
rect 12182 22120 12188 22172
rect 55062 22120 55068 22172
rect 55120 22120 55126 22172
rect 12124 21880 12130 21932
rect 12182 21880 12188 21932
rect 55062 21880 55068 21932
rect 55120 21880 55126 21932
rect 12124 21330 12130 21382
rect 12182 21330 12188 21382
rect 55062 21330 55068 21382
rect 55120 21330 55126 21382
rect 12124 21090 12130 21142
rect 12182 21090 12188 21142
rect 55062 21090 55068 21142
rect 55120 21090 55126 21142
rect 12124 20540 12130 20592
rect 12182 20540 12188 20592
rect 55062 20540 55068 20592
rect 55120 20540 55126 20592
rect 12124 20300 12130 20352
rect 12182 20300 12188 20352
rect 55062 20300 55068 20352
rect 55120 20300 55126 20352
rect 12124 19750 12130 19802
rect 12182 19750 12188 19802
rect 55062 19750 55068 19802
rect 55120 19750 55126 19802
rect 12124 19510 12130 19562
rect 12182 19510 12188 19562
rect 55062 19510 55068 19562
rect 55120 19510 55126 19562
rect 12124 18960 12130 19012
rect 12182 18960 12188 19012
rect 55062 18960 55068 19012
rect 55120 18960 55126 19012
rect 12124 18720 12130 18772
rect 12182 18720 12188 18772
rect 55062 18720 55068 18772
rect 55120 18720 55126 18772
rect 12124 18170 12130 18222
rect 12182 18170 12188 18222
rect 55062 18170 55068 18222
rect 55120 18170 55126 18222
rect 19 10176 47 18076
rect 99 10176 127 18076
rect 179 10176 207 18076
rect 259 10176 287 18076
rect 339 10176 367 18076
rect 419 10176 447 18076
rect 499 10176 527 18076
rect 12124 17930 12130 17982
rect 12182 17930 12188 17982
rect 55062 17930 55068 17982
rect 55120 17930 55126 17982
rect 12124 17380 12130 17432
rect 12182 17380 12188 17432
rect 55062 17380 55068 17432
rect 55120 17380 55126 17432
rect 12124 17140 12130 17192
rect 12182 17140 12188 17192
rect 55062 17140 55068 17192
rect 55120 17140 55126 17192
rect 12124 16590 12130 16642
rect 12182 16590 12188 16642
rect 55062 16590 55068 16642
rect 55120 16590 55126 16642
rect 12124 16350 12130 16402
rect 12182 16350 12188 16402
rect 55062 16350 55068 16402
rect 55120 16350 55126 16402
rect 12124 15800 12130 15852
rect 12182 15800 12188 15852
rect 55062 15800 55068 15852
rect 55120 15800 55126 15852
rect 12124 15560 12130 15612
rect 12182 15560 12188 15612
rect 55062 15560 55068 15612
rect 55120 15560 55126 15612
rect 12124 15010 12130 15062
rect 12182 15010 12188 15062
rect 55062 15010 55068 15062
rect 55120 15010 55126 15062
rect 12124 14770 12130 14822
rect 12182 14770 12188 14822
rect 55062 14770 55068 14822
rect 55120 14770 55126 14822
rect 12124 14220 12130 14272
rect 12182 14220 12188 14272
rect 55062 14220 55068 14272
rect 55120 14220 55126 14272
rect 12124 13980 12130 14032
rect 12182 13980 12188 14032
rect 55062 13980 55068 14032
rect 55120 13980 55126 14032
rect 12124 13430 12130 13482
rect 12182 13430 12188 13482
rect 55062 13430 55068 13482
rect 55120 13430 55126 13482
rect 12124 13190 12130 13242
rect 12182 13190 12188 13242
rect 55062 13190 55068 13242
rect 55120 13190 55126 13242
rect 12124 12640 12130 12692
rect 12182 12640 12188 12692
rect 55062 12640 55068 12692
rect 55120 12640 55126 12692
rect 12124 12400 12130 12452
rect 12182 12400 12188 12452
rect 55062 12400 55068 12452
rect 55120 12400 55126 12452
rect 12124 11850 12130 11902
rect 12182 11850 12188 11902
rect 55062 11850 55068 11902
rect 55120 11850 55126 11902
rect 12124 11610 12130 11662
rect 12182 11610 12188 11662
rect 55062 11610 55068 11662
rect 55120 11610 55126 11662
rect 12124 11060 12130 11112
rect 12182 11060 12188 11112
rect 55062 11060 55068 11112
rect 55120 11060 55126 11112
rect 12124 10820 12130 10872
rect 12182 10820 12188 10872
rect 55062 10820 55068 10872
rect 55120 10820 55126 10872
rect 12124 10270 12130 10322
rect 12182 10270 12188 10322
rect 55062 10270 55068 10322
rect 55120 10270 55126 10322
rect 66723 10176 66751 18076
rect 66803 10176 66831 18076
rect 66883 10176 66911 18076
rect 66963 10176 66991 18076
rect 67043 10176 67071 18076
rect 67123 10176 67151 18076
rect 67203 10176 67231 18076
rect 12124 10030 12130 10082
rect 12182 10030 12188 10082
rect 13475 9274 13503 9386
rect 13099 9246 13503 9274
rect 13547 9274 13575 9386
rect 13739 9274 13767 9386
rect 13547 9246 13591 9274
rect 13099 9134 13127 9246
rect 13563 9134 13591 9246
rect 13723 9246 13767 9274
rect 13811 9274 13839 9386
rect 14723 9274 14751 9386
rect 13811 9246 14215 9274
rect 13723 9134 13751 9246
rect 14187 9134 14215 9246
rect 14347 9246 14751 9274
rect 14795 9274 14823 9386
rect 14987 9274 15015 9386
rect 14795 9246 14839 9274
rect 14347 9134 14375 9246
rect 14811 9134 14839 9246
rect 14971 9246 15015 9274
rect 15059 9274 15087 9386
rect 15971 9274 15999 9386
rect 15059 9246 15463 9274
rect 14971 9134 14999 9246
rect 15435 9134 15463 9246
rect 15595 9246 15999 9274
rect 16043 9274 16071 9386
rect 16235 9274 16263 9386
rect 16043 9246 16087 9274
rect 15595 9134 15623 9246
rect 16059 9134 16087 9246
rect 16219 9246 16263 9274
rect 16307 9274 16335 9386
rect 17219 9274 17247 9386
rect 16307 9246 16711 9274
rect 16219 9134 16247 9246
rect 16683 9134 16711 9246
rect 16843 9246 17247 9274
rect 17291 9274 17319 9386
rect 17483 9274 17511 9386
rect 17291 9246 17335 9274
rect 16843 9134 16871 9246
rect 17307 9134 17335 9246
rect 17467 9246 17511 9274
rect 17555 9274 17583 9386
rect 18467 9274 18495 9386
rect 17555 9246 17959 9274
rect 17467 9134 17495 9246
rect 17931 9134 17959 9246
rect 18091 9246 18495 9274
rect 18539 9274 18567 9386
rect 18731 9274 18759 9386
rect 18539 9246 18583 9274
rect 18091 9134 18119 9246
rect 18555 9134 18583 9246
rect 18715 9246 18759 9274
rect 18803 9274 18831 9386
rect 19715 9274 19743 9386
rect 18803 9246 19207 9274
rect 18715 9134 18743 9246
rect 19179 9134 19207 9246
rect 19339 9246 19743 9274
rect 19787 9274 19815 9386
rect 19979 9274 20007 9386
rect 19787 9246 19831 9274
rect 19339 9134 19367 9246
rect 19803 9134 19831 9246
rect 19963 9246 20007 9274
rect 20051 9274 20079 9386
rect 20963 9274 20991 9386
rect 20051 9246 20455 9274
rect 19963 9134 19991 9246
rect 20427 9134 20455 9246
rect 20587 9246 20991 9274
rect 21035 9274 21063 9386
rect 21227 9274 21255 9386
rect 21035 9246 21079 9274
rect 20587 9134 20615 9246
rect 21051 9134 21079 9246
rect 21211 9246 21255 9274
rect 21299 9274 21327 9386
rect 22211 9274 22239 9386
rect 21299 9246 21703 9274
rect 21211 9134 21239 9246
rect 21675 9134 21703 9246
rect 21835 9246 22239 9274
rect 22283 9274 22311 9386
rect 22475 9274 22503 9386
rect 22283 9246 22327 9274
rect 21835 9134 21863 9246
rect 22299 9134 22327 9246
rect 22459 9246 22503 9274
rect 22547 9274 22575 9386
rect 23459 9274 23487 9386
rect 22547 9246 22951 9274
rect 22459 9134 22487 9246
rect 22923 9134 22951 9246
rect 23083 9246 23487 9274
rect 23531 9274 23559 9386
rect 23723 9274 23751 9386
rect 23531 9246 23575 9274
rect 23083 9134 23111 9246
rect 23547 9134 23575 9246
rect 23707 9246 23751 9274
rect 23795 9274 23823 9386
rect 24707 9274 24735 9386
rect 23795 9246 24199 9274
rect 23707 9134 23735 9246
rect 24171 9134 24199 9246
rect 24331 9246 24735 9274
rect 24779 9274 24807 9386
rect 24971 9274 24999 9386
rect 24779 9246 24823 9274
rect 24331 9134 24359 9246
rect 24795 9134 24823 9246
rect 24955 9246 24999 9274
rect 25043 9274 25071 9386
rect 25955 9274 25983 9386
rect 25043 9246 25447 9274
rect 24955 9134 24983 9246
rect 25419 9134 25447 9246
rect 25579 9246 25983 9274
rect 26027 9274 26055 9386
rect 26219 9274 26247 9386
rect 26027 9246 26071 9274
rect 25579 9134 25607 9246
rect 26043 9134 26071 9246
rect 26203 9246 26247 9274
rect 26291 9274 26319 9386
rect 27203 9274 27231 9386
rect 26291 9246 26695 9274
rect 26203 9134 26231 9246
rect 26667 9134 26695 9246
rect 26827 9246 27231 9274
rect 27275 9274 27303 9386
rect 27467 9274 27495 9386
rect 27275 9246 27319 9274
rect 26827 9134 26855 9246
rect 27291 9134 27319 9246
rect 27451 9246 27495 9274
rect 27539 9274 27567 9386
rect 28451 9274 28479 9386
rect 27539 9246 27943 9274
rect 27451 9134 27479 9246
rect 27915 9134 27943 9246
rect 28075 9246 28479 9274
rect 28523 9274 28551 9386
rect 28715 9274 28743 9386
rect 28523 9246 28567 9274
rect 28075 9134 28103 9246
rect 28539 9134 28567 9246
rect 28699 9246 28743 9274
rect 28787 9274 28815 9386
rect 29699 9274 29727 9386
rect 28787 9246 29191 9274
rect 28699 9134 28727 9246
rect 29163 9134 29191 9246
rect 29323 9246 29727 9274
rect 29771 9274 29799 9386
rect 29963 9274 29991 9386
rect 29771 9246 29815 9274
rect 29323 9134 29351 9246
rect 29787 9134 29815 9246
rect 29947 9246 29991 9274
rect 30035 9274 30063 9386
rect 30947 9274 30975 9386
rect 30035 9246 30439 9274
rect 29947 9134 29975 9246
rect 30411 9134 30439 9246
rect 30571 9246 30975 9274
rect 31019 9274 31047 9386
rect 31211 9274 31239 9386
rect 31019 9246 31063 9274
rect 30571 9134 30599 9246
rect 31035 9134 31063 9246
rect 31195 9246 31239 9274
rect 31283 9274 31311 9386
rect 32195 9274 32223 9386
rect 31283 9246 31687 9274
rect 31195 9134 31223 9246
rect 31659 9134 31687 9246
rect 31819 9246 32223 9274
rect 32267 9274 32295 9386
rect 32459 9274 32487 9386
rect 32267 9246 32311 9274
rect 31819 9134 31847 9246
rect 32283 9134 32311 9246
rect 32443 9246 32487 9274
rect 32531 9274 32559 9386
rect 33443 9274 33471 9386
rect 32531 9246 32935 9274
rect 32443 9134 32471 9246
rect 32907 9134 32935 9246
rect 33067 9246 33471 9274
rect 33515 9274 33543 9386
rect 33707 9274 33735 9386
rect 33515 9246 33559 9274
rect 33067 9134 33095 9246
rect 33531 9134 33559 9246
rect 33691 9246 33735 9274
rect 33779 9274 33807 9386
rect 34691 9274 34719 9386
rect 33779 9246 34183 9274
rect 33691 9134 33719 9246
rect 34155 9134 34183 9246
rect 34315 9246 34719 9274
rect 34763 9274 34791 9386
rect 34955 9274 34983 9386
rect 34763 9246 34807 9274
rect 34315 9134 34343 9246
rect 34779 9134 34807 9246
rect 34939 9246 34983 9274
rect 35027 9274 35055 9386
rect 35939 9274 35967 9386
rect 35027 9246 35431 9274
rect 34939 9134 34967 9246
rect 35403 9134 35431 9246
rect 35563 9246 35967 9274
rect 36011 9274 36039 9386
rect 36203 9274 36231 9386
rect 36011 9246 36055 9274
rect 35563 9134 35591 9246
rect 36027 9134 36055 9246
rect 36187 9246 36231 9274
rect 36275 9274 36303 9386
rect 37187 9274 37215 9386
rect 36275 9246 36679 9274
rect 36187 9134 36215 9246
rect 36651 9134 36679 9246
rect 36811 9246 37215 9274
rect 37259 9274 37287 9386
rect 37451 9274 37479 9386
rect 37259 9246 37303 9274
rect 36811 9134 36839 9246
rect 37275 9134 37303 9246
rect 37435 9246 37479 9274
rect 37523 9274 37551 9386
rect 38435 9274 38463 9386
rect 37523 9246 37927 9274
rect 37435 9134 37463 9246
rect 37899 9134 37927 9246
rect 38059 9246 38463 9274
rect 38507 9274 38535 9386
rect 38699 9274 38727 9386
rect 38507 9246 38551 9274
rect 38059 9134 38087 9246
rect 38523 9134 38551 9246
rect 38683 9246 38727 9274
rect 38771 9274 38799 9386
rect 39683 9274 39711 9386
rect 38771 9246 39175 9274
rect 38683 9134 38711 9246
rect 39147 9134 39175 9246
rect 39307 9246 39711 9274
rect 39755 9274 39783 9386
rect 39947 9274 39975 9386
rect 39755 9246 39799 9274
rect 39307 9134 39335 9246
rect 39771 9134 39799 9246
rect 39931 9246 39975 9274
rect 40019 9274 40047 9386
rect 40931 9274 40959 9386
rect 40019 9246 40423 9274
rect 39931 9134 39959 9246
rect 40395 9134 40423 9246
rect 40555 9246 40959 9274
rect 41003 9274 41031 9386
rect 41195 9274 41223 9386
rect 41003 9246 41047 9274
rect 40555 9134 40583 9246
rect 41019 9134 41047 9246
rect 41179 9246 41223 9274
rect 41267 9274 41295 9386
rect 42179 9274 42207 9386
rect 41267 9246 41671 9274
rect 41179 9134 41207 9246
rect 41643 9134 41671 9246
rect 41803 9246 42207 9274
rect 42251 9274 42279 9386
rect 42443 9274 42471 9386
rect 42251 9246 42295 9274
rect 41803 9134 41831 9246
rect 42267 9134 42295 9246
rect 42427 9246 42471 9274
rect 42515 9274 42543 9386
rect 43427 9274 43455 9386
rect 42515 9246 42919 9274
rect 42427 9134 42455 9246
rect 42891 9134 42919 9246
rect 43051 9246 43455 9274
rect 43499 9274 43527 9386
rect 43691 9274 43719 9386
rect 43499 9246 43543 9274
rect 43051 9134 43079 9246
rect 43515 9134 43543 9246
rect 43675 9246 43719 9274
rect 43763 9274 43791 9386
rect 44675 9274 44703 9386
rect 43763 9246 44167 9274
rect 43675 9134 43703 9246
rect 44139 9134 44167 9246
rect 44299 9246 44703 9274
rect 44747 9274 44775 9386
rect 44939 9274 44967 9386
rect 44747 9246 44791 9274
rect 44299 9134 44327 9246
rect 44763 9134 44791 9246
rect 44923 9246 44967 9274
rect 45011 9274 45039 9386
rect 45923 9274 45951 9386
rect 45011 9246 45415 9274
rect 44923 9134 44951 9246
rect 45387 9134 45415 9246
rect 45547 9246 45951 9274
rect 45995 9274 46023 9386
rect 46187 9274 46215 9386
rect 45995 9246 46039 9274
rect 45547 9134 45575 9246
rect 46011 9134 46039 9246
rect 46171 9246 46215 9274
rect 46259 9274 46287 9386
rect 47171 9274 47199 9386
rect 46259 9246 46663 9274
rect 46171 9134 46199 9246
rect 46635 9134 46663 9246
rect 46795 9246 47199 9274
rect 47243 9274 47271 9386
rect 47435 9274 47463 9386
rect 47243 9246 47287 9274
rect 46795 9134 46823 9246
rect 47259 9134 47287 9246
rect 47419 9246 47463 9274
rect 47507 9274 47535 9386
rect 48419 9274 48447 9386
rect 47507 9246 47911 9274
rect 47419 9134 47447 9246
rect 47883 9134 47911 9246
rect 48043 9246 48447 9274
rect 48491 9274 48519 9386
rect 48683 9274 48711 9386
rect 48491 9246 48535 9274
rect 48043 9134 48071 9246
rect 48507 9134 48535 9246
rect 48667 9246 48711 9274
rect 48755 9274 48783 9386
rect 49667 9274 49695 9386
rect 48755 9246 49159 9274
rect 48667 9134 48695 9246
rect 49131 9134 49159 9246
rect 49291 9246 49695 9274
rect 49739 9274 49767 9386
rect 49931 9274 49959 9386
rect 49739 9246 49783 9274
rect 49291 9134 49319 9246
rect 49755 9134 49783 9246
rect 49915 9246 49959 9274
rect 50003 9274 50031 9386
rect 50915 9274 50943 9386
rect 50003 9246 50407 9274
rect 49915 9134 49943 9246
rect 50379 9134 50407 9246
rect 50539 9246 50943 9274
rect 50987 9274 51015 9386
rect 51179 9274 51207 9386
rect 50987 9246 51031 9274
rect 50539 9134 50567 9246
rect 51003 9134 51031 9246
rect 51163 9246 51207 9274
rect 51251 9274 51279 9386
rect 52163 9274 52191 9386
rect 51251 9246 51655 9274
rect 51163 9134 51191 9246
rect 51627 9134 51655 9246
rect 51787 9246 52191 9274
rect 52235 9274 52263 9386
rect 52427 9274 52455 9386
rect 52235 9246 52279 9274
rect 51787 9134 51815 9246
rect 52251 9134 52279 9246
rect 52411 9246 52455 9274
rect 52499 9274 52527 9386
rect 53411 9274 53439 9386
rect 52499 9246 52903 9274
rect 52411 9134 52439 9246
rect 52875 9134 52903 9246
rect 53035 9246 53439 9274
rect 53483 9274 53511 9386
rect 53483 9246 53527 9274
rect 53035 9134 53063 9246
rect 53499 9134 53527 9246
rect 13563 8282 13591 8380
rect 13545 8230 13551 8282
rect 13603 8230 13609 8282
rect 6725 7609 6731 7661
rect 6783 7609 6789 7661
rect 7124 6902 7130 6954
rect 7182 6902 7188 6954
rect 6725 6195 6731 6247
rect 6783 6195 6789 6247
rect 7124 5488 7130 5540
rect 7182 5488 7188 5540
rect 6725 4781 6731 4833
rect 6783 4781 6789 4833
rect 13761 3684 13807 3938
rect 15009 3684 15055 3938
rect 16257 3684 16303 3938
rect 17505 3684 17551 3938
rect 18753 3684 18799 3938
rect 20001 3684 20047 3938
rect 21249 3684 21295 3938
rect 22497 3684 22543 3938
rect 23745 3684 23791 3938
rect 24993 3684 25039 3938
rect 26241 3684 26287 3938
rect 27489 3684 27535 3938
rect 28737 3684 28783 3938
rect 29985 3684 30031 3938
rect 31233 3684 31279 3938
rect 32481 3684 32527 3938
rect 33729 3684 33775 3938
rect 34977 3684 35023 3938
rect 36225 3684 36271 3938
rect 37473 3684 37519 3938
rect 38721 3684 38767 3938
rect 39969 3684 40015 3938
rect 41217 3684 41263 3938
rect 42465 3684 42511 3938
rect 43713 3684 43759 3938
rect 44961 3684 45007 3938
rect 46209 3684 46255 3938
rect 47457 3684 47503 3938
rect 48705 3684 48751 3938
rect 49953 3684 49999 3938
rect 51201 3684 51247 3938
rect 52449 3684 52495 3938
rect 13912 1425 13972 1481
rect 15160 1425 15220 1481
rect 16408 1425 16468 1481
rect 17656 1425 17716 1481
rect 18904 1425 18964 1481
rect 20152 1425 20212 1481
rect 21400 1425 21460 1481
rect 22648 1425 22708 1481
rect 23896 1425 23956 1481
rect 25144 1425 25204 1481
rect 26392 1425 26452 1481
rect 27640 1425 27700 1481
rect 28888 1425 28948 1481
rect 30136 1425 30196 1481
rect 31384 1425 31444 1481
rect 32632 1425 32692 1481
rect 33880 1425 33940 1481
rect 35128 1425 35188 1481
rect 36376 1425 36436 1481
rect 37624 1425 37684 1481
rect 38872 1425 38932 1481
rect 40120 1425 40180 1481
rect 41368 1425 41428 1481
rect 42616 1425 42676 1481
rect 43864 1425 43924 1481
rect 45112 1425 45172 1481
rect 46360 1425 46420 1481
rect 47608 1425 47668 1481
rect 48856 1425 48916 1481
rect 50104 1425 50164 1481
rect 51352 1425 51412 1481
rect 52600 1425 52660 1481
<< via1 >>
rect 60343 66122 60395 66131
rect 60343 66088 60352 66122
rect 60352 66088 60386 66122
rect 60386 66088 60395 66122
rect 60343 66079 60395 66088
rect 59944 65415 59996 65424
rect 59944 65381 59953 65415
rect 59953 65381 59987 65415
rect 59987 65381 59996 65415
rect 59944 65372 59996 65381
rect 60343 64708 60395 64717
rect 60343 64674 60352 64708
rect 60352 64674 60386 64708
rect 60386 64674 60395 64708
rect 60343 64665 60395 64674
rect 59944 64001 59996 64010
rect 59944 63967 59953 64001
rect 59953 63967 59987 64001
rect 59987 63967 59996 64001
rect 59944 63958 59996 63967
rect 60343 63294 60395 63303
rect 60343 63260 60352 63294
rect 60352 63260 60386 63294
rect 60386 63260 60395 63294
rect 60343 63251 60395 63260
rect 53647 62630 53699 62682
rect 55068 60873 55120 60882
rect 55068 60839 55077 60873
rect 55077 60839 55111 60873
rect 55111 60839 55120 60873
rect 55068 60830 55120 60839
rect 12130 60633 12182 60642
rect 12130 60599 12139 60633
rect 12139 60599 12173 60633
rect 12173 60599 12182 60633
rect 12130 60590 12182 60599
rect 55068 60633 55120 60642
rect 55068 60599 55077 60633
rect 55077 60599 55111 60633
rect 55111 60599 55120 60633
rect 55068 60590 55120 60599
rect 12130 60083 12182 60092
rect 12130 60049 12139 60083
rect 12139 60049 12173 60083
rect 12173 60049 12182 60083
rect 12130 60040 12182 60049
rect 55068 60083 55120 60092
rect 55068 60049 55077 60083
rect 55077 60049 55111 60083
rect 55111 60049 55120 60083
rect 55068 60040 55120 60049
rect 12130 59843 12182 59852
rect 12130 59809 12139 59843
rect 12139 59809 12173 59843
rect 12173 59809 12182 59843
rect 12130 59800 12182 59809
rect 55068 59843 55120 59852
rect 55068 59809 55077 59843
rect 55077 59809 55111 59843
rect 55111 59809 55120 59843
rect 55068 59800 55120 59809
rect 12130 59293 12182 59302
rect 12130 59259 12139 59293
rect 12139 59259 12173 59293
rect 12173 59259 12182 59293
rect 12130 59250 12182 59259
rect 55068 59293 55120 59302
rect 55068 59259 55077 59293
rect 55077 59259 55111 59293
rect 55111 59259 55120 59293
rect 55068 59250 55120 59259
rect 12130 59053 12182 59062
rect 12130 59019 12139 59053
rect 12139 59019 12173 59053
rect 12173 59019 12182 59053
rect 12130 59010 12182 59019
rect 55068 59053 55120 59062
rect 55068 59019 55077 59053
rect 55077 59019 55111 59053
rect 55111 59019 55120 59053
rect 55068 59010 55120 59019
rect 12130 58503 12182 58512
rect 12130 58469 12139 58503
rect 12139 58469 12173 58503
rect 12173 58469 12182 58503
rect 12130 58460 12182 58469
rect 55068 58503 55120 58512
rect 55068 58469 55077 58503
rect 55077 58469 55111 58503
rect 55111 58469 55120 58503
rect 55068 58460 55120 58469
rect 12130 58263 12182 58272
rect 12130 58229 12139 58263
rect 12139 58229 12173 58263
rect 12173 58229 12182 58263
rect 12130 58220 12182 58229
rect 55068 58263 55120 58272
rect 55068 58229 55077 58263
rect 55077 58229 55111 58263
rect 55111 58229 55120 58263
rect 55068 58220 55120 58229
rect 12130 57713 12182 57722
rect 12130 57679 12139 57713
rect 12139 57679 12173 57713
rect 12173 57679 12182 57713
rect 12130 57670 12182 57679
rect 55068 57713 55120 57722
rect 55068 57679 55077 57713
rect 55077 57679 55111 57713
rect 55111 57679 55120 57713
rect 55068 57670 55120 57679
rect 12130 57473 12182 57482
rect 12130 57439 12139 57473
rect 12139 57439 12173 57473
rect 12173 57439 12182 57473
rect 12130 57430 12182 57439
rect 55068 57473 55120 57482
rect 55068 57439 55077 57473
rect 55077 57439 55111 57473
rect 55111 57439 55120 57473
rect 55068 57430 55120 57439
rect 12130 56923 12182 56932
rect 12130 56889 12139 56923
rect 12139 56889 12173 56923
rect 12173 56889 12182 56923
rect 12130 56880 12182 56889
rect 55068 56923 55120 56932
rect 55068 56889 55077 56923
rect 55077 56889 55111 56923
rect 55111 56889 55120 56923
rect 55068 56880 55120 56889
rect 12130 56683 12182 56692
rect 12130 56649 12139 56683
rect 12139 56649 12173 56683
rect 12173 56649 12182 56683
rect 12130 56640 12182 56649
rect 55068 56683 55120 56692
rect 55068 56649 55077 56683
rect 55077 56649 55111 56683
rect 55111 56649 55120 56683
rect 55068 56640 55120 56649
rect 12130 56133 12182 56142
rect 12130 56099 12139 56133
rect 12139 56099 12173 56133
rect 12173 56099 12182 56133
rect 12130 56090 12182 56099
rect 55068 56133 55120 56142
rect 55068 56099 55077 56133
rect 55077 56099 55111 56133
rect 55111 56099 55120 56133
rect 55068 56090 55120 56099
rect 12130 55893 12182 55902
rect 12130 55859 12139 55893
rect 12139 55859 12173 55893
rect 12173 55859 12182 55893
rect 12130 55850 12182 55859
rect 55068 55893 55120 55902
rect 55068 55859 55077 55893
rect 55077 55859 55111 55893
rect 55111 55859 55120 55893
rect 55068 55850 55120 55859
rect 12130 55343 12182 55352
rect 12130 55309 12139 55343
rect 12139 55309 12173 55343
rect 12173 55309 12182 55343
rect 12130 55300 12182 55309
rect 55068 55343 55120 55352
rect 55068 55309 55077 55343
rect 55077 55309 55111 55343
rect 55111 55309 55120 55343
rect 55068 55300 55120 55309
rect 12130 55103 12182 55112
rect 12130 55069 12139 55103
rect 12139 55069 12173 55103
rect 12173 55069 12182 55103
rect 12130 55060 12182 55069
rect 55068 55103 55120 55112
rect 55068 55069 55077 55103
rect 55077 55069 55111 55103
rect 55111 55069 55120 55103
rect 55068 55060 55120 55069
rect 12130 54553 12182 54562
rect 12130 54519 12139 54553
rect 12139 54519 12173 54553
rect 12173 54519 12182 54553
rect 12130 54510 12182 54519
rect 55068 54553 55120 54562
rect 55068 54519 55077 54553
rect 55077 54519 55111 54553
rect 55111 54519 55120 54553
rect 55068 54510 55120 54519
rect 12130 54313 12182 54322
rect 12130 54279 12139 54313
rect 12139 54279 12173 54313
rect 12173 54279 12182 54313
rect 12130 54270 12182 54279
rect 55068 54313 55120 54322
rect 55068 54279 55077 54313
rect 55077 54279 55111 54313
rect 55111 54279 55120 54313
rect 55068 54270 55120 54279
rect 12130 53763 12182 53772
rect 12130 53729 12139 53763
rect 12139 53729 12173 53763
rect 12173 53729 12182 53763
rect 12130 53720 12182 53729
rect 55068 53763 55120 53772
rect 55068 53729 55077 53763
rect 55077 53729 55111 53763
rect 55111 53729 55120 53763
rect 55068 53720 55120 53729
rect 12130 53523 12182 53532
rect 12130 53489 12139 53523
rect 12139 53489 12173 53523
rect 12173 53489 12182 53523
rect 12130 53480 12182 53489
rect 55068 53523 55120 53532
rect 55068 53489 55077 53523
rect 55077 53489 55111 53523
rect 55111 53489 55120 53523
rect 55068 53480 55120 53489
rect 12130 52973 12182 52982
rect 12130 52939 12139 52973
rect 12139 52939 12173 52973
rect 12173 52939 12182 52973
rect 12130 52930 12182 52939
rect 55068 52973 55120 52982
rect 55068 52939 55077 52973
rect 55077 52939 55111 52973
rect 55111 52939 55120 52973
rect 55068 52930 55120 52939
rect 12130 52733 12182 52742
rect 12130 52699 12139 52733
rect 12139 52699 12173 52733
rect 12173 52699 12182 52733
rect 12130 52690 12182 52699
rect 55068 52733 55120 52742
rect 55068 52699 55077 52733
rect 55077 52699 55111 52733
rect 55111 52699 55120 52733
rect 55068 52690 55120 52699
rect 12130 52183 12182 52192
rect 12130 52149 12139 52183
rect 12139 52149 12173 52183
rect 12173 52149 12182 52183
rect 12130 52140 12182 52149
rect 55068 52183 55120 52192
rect 55068 52149 55077 52183
rect 55077 52149 55111 52183
rect 55111 52149 55120 52183
rect 55068 52140 55120 52149
rect 12130 51943 12182 51952
rect 12130 51909 12139 51943
rect 12139 51909 12173 51943
rect 12173 51909 12182 51943
rect 12130 51900 12182 51909
rect 55068 51943 55120 51952
rect 55068 51909 55077 51943
rect 55077 51909 55111 51943
rect 55111 51909 55120 51943
rect 55068 51900 55120 51909
rect 12130 51393 12182 51402
rect 12130 51359 12139 51393
rect 12139 51359 12173 51393
rect 12173 51359 12182 51393
rect 12130 51350 12182 51359
rect 55068 51393 55120 51402
rect 55068 51359 55077 51393
rect 55077 51359 55111 51393
rect 55111 51359 55120 51393
rect 55068 51350 55120 51359
rect 12130 51153 12182 51162
rect 12130 51119 12139 51153
rect 12139 51119 12173 51153
rect 12173 51119 12182 51153
rect 12130 51110 12182 51119
rect 55068 51153 55120 51162
rect 55068 51119 55077 51153
rect 55077 51119 55111 51153
rect 55111 51119 55120 51153
rect 55068 51110 55120 51119
rect 12130 50603 12182 50612
rect 12130 50569 12139 50603
rect 12139 50569 12173 50603
rect 12173 50569 12182 50603
rect 12130 50560 12182 50569
rect 55068 50603 55120 50612
rect 55068 50569 55077 50603
rect 55077 50569 55111 50603
rect 55111 50569 55120 50603
rect 55068 50560 55120 50569
rect 12130 50363 12182 50372
rect 12130 50329 12139 50363
rect 12139 50329 12173 50363
rect 12173 50329 12182 50363
rect 12130 50320 12182 50329
rect 55068 50363 55120 50372
rect 55068 50329 55077 50363
rect 55077 50329 55111 50363
rect 55111 50329 55120 50363
rect 55068 50320 55120 50329
rect 12130 49813 12182 49822
rect 12130 49779 12139 49813
rect 12139 49779 12173 49813
rect 12173 49779 12182 49813
rect 12130 49770 12182 49779
rect 55068 49813 55120 49822
rect 55068 49779 55077 49813
rect 55077 49779 55111 49813
rect 55111 49779 55120 49813
rect 55068 49770 55120 49779
rect 12130 49573 12182 49582
rect 12130 49539 12139 49573
rect 12139 49539 12173 49573
rect 12173 49539 12182 49573
rect 12130 49530 12182 49539
rect 55068 49573 55120 49582
rect 55068 49539 55077 49573
rect 55077 49539 55111 49573
rect 55111 49539 55120 49573
rect 55068 49530 55120 49539
rect 12130 49023 12182 49032
rect 12130 48989 12139 49023
rect 12139 48989 12173 49023
rect 12173 48989 12182 49023
rect 12130 48980 12182 48989
rect 55068 49023 55120 49032
rect 55068 48989 55077 49023
rect 55077 48989 55111 49023
rect 55111 48989 55120 49023
rect 55068 48980 55120 48989
rect 12130 48783 12182 48792
rect 12130 48749 12139 48783
rect 12139 48749 12173 48783
rect 12173 48749 12182 48783
rect 12130 48740 12182 48749
rect 55068 48783 55120 48792
rect 55068 48749 55077 48783
rect 55077 48749 55111 48783
rect 55111 48749 55120 48783
rect 55068 48740 55120 48749
rect 12130 48233 12182 48242
rect 12130 48199 12139 48233
rect 12139 48199 12173 48233
rect 12173 48199 12182 48233
rect 12130 48190 12182 48199
rect 55068 48233 55120 48242
rect 55068 48199 55077 48233
rect 55077 48199 55111 48233
rect 55111 48199 55120 48233
rect 55068 48190 55120 48199
rect 12130 47993 12182 48002
rect 12130 47959 12139 47993
rect 12139 47959 12173 47993
rect 12173 47959 12182 47993
rect 12130 47950 12182 47959
rect 55068 47993 55120 48002
rect 55068 47959 55077 47993
rect 55077 47959 55111 47993
rect 55111 47959 55120 47993
rect 55068 47950 55120 47959
rect 12130 47443 12182 47452
rect 12130 47409 12139 47443
rect 12139 47409 12173 47443
rect 12173 47409 12182 47443
rect 12130 47400 12182 47409
rect 55068 47443 55120 47452
rect 55068 47409 55077 47443
rect 55077 47409 55111 47443
rect 55111 47409 55120 47443
rect 55068 47400 55120 47409
rect 12130 47203 12182 47212
rect 12130 47169 12139 47203
rect 12139 47169 12173 47203
rect 12173 47169 12182 47203
rect 12130 47160 12182 47169
rect 55068 47203 55120 47212
rect 55068 47169 55077 47203
rect 55077 47169 55111 47203
rect 55111 47169 55120 47203
rect 55068 47160 55120 47169
rect 12130 46653 12182 46662
rect 12130 46619 12139 46653
rect 12139 46619 12173 46653
rect 12173 46619 12182 46653
rect 12130 46610 12182 46619
rect 55068 46653 55120 46662
rect 55068 46619 55077 46653
rect 55077 46619 55111 46653
rect 55111 46619 55120 46653
rect 55068 46610 55120 46619
rect 12130 46413 12182 46422
rect 12130 46379 12139 46413
rect 12139 46379 12173 46413
rect 12173 46379 12182 46413
rect 12130 46370 12182 46379
rect 55068 46413 55120 46422
rect 55068 46379 55077 46413
rect 55077 46379 55111 46413
rect 55111 46379 55120 46413
rect 55068 46370 55120 46379
rect 12130 45863 12182 45872
rect 12130 45829 12139 45863
rect 12139 45829 12173 45863
rect 12173 45829 12182 45863
rect 12130 45820 12182 45829
rect 55068 45863 55120 45872
rect 55068 45829 55077 45863
rect 55077 45829 55111 45863
rect 55111 45829 55120 45863
rect 55068 45820 55120 45829
rect 12130 45623 12182 45632
rect 12130 45589 12139 45623
rect 12139 45589 12173 45623
rect 12173 45589 12182 45623
rect 12130 45580 12182 45589
rect 55068 45623 55120 45632
rect 55068 45589 55077 45623
rect 55077 45589 55111 45623
rect 55111 45589 55120 45623
rect 55068 45580 55120 45589
rect 12130 45073 12182 45082
rect 12130 45039 12139 45073
rect 12139 45039 12173 45073
rect 12173 45039 12182 45073
rect 12130 45030 12182 45039
rect 55068 45073 55120 45082
rect 55068 45039 55077 45073
rect 55077 45039 55111 45073
rect 55111 45039 55120 45073
rect 55068 45030 55120 45039
rect 12130 44833 12182 44842
rect 12130 44799 12139 44833
rect 12139 44799 12173 44833
rect 12173 44799 12182 44833
rect 12130 44790 12182 44799
rect 55068 44833 55120 44842
rect 55068 44799 55077 44833
rect 55077 44799 55111 44833
rect 55111 44799 55120 44833
rect 55068 44790 55120 44799
rect 12130 44283 12182 44292
rect 12130 44249 12139 44283
rect 12139 44249 12173 44283
rect 12173 44249 12182 44283
rect 12130 44240 12182 44249
rect 55068 44283 55120 44292
rect 55068 44249 55077 44283
rect 55077 44249 55111 44283
rect 55111 44249 55120 44283
rect 55068 44240 55120 44249
rect 12130 44043 12182 44052
rect 12130 44009 12139 44043
rect 12139 44009 12173 44043
rect 12173 44009 12182 44043
rect 12130 44000 12182 44009
rect 55068 44043 55120 44052
rect 55068 44009 55077 44043
rect 55077 44009 55111 44043
rect 55111 44009 55120 44043
rect 55068 44000 55120 44009
rect 12130 43493 12182 43502
rect 12130 43459 12139 43493
rect 12139 43459 12173 43493
rect 12173 43459 12182 43493
rect 12130 43450 12182 43459
rect 55068 43493 55120 43502
rect 55068 43459 55077 43493
rect 55077 43459 55111 43493
rect 55111 43459 55120 43493
rect 55068 43450 55120 43459
rect 12130 43253 12182 43262
rect 12130 43219 12139 43253
rect 12139 43219 12173 43253
rect 12173 43219 12182 43253
rect 12130 43210 12182 43219
rect 55068 43253 55120 43262
rect 55068 43219 55077 43253
rect 55077 43219 55111 43253
rect 55111 43219 55120 43253
rect 55068 43210 55120 43219
rect 12130 42703 12182 42712
rect 12130 42669 12139 42703
rect 12139 42669 12173 42703
rect 12173 42669 12182 42703
rect 12130 42660 12182 42669
rect 55068 42703 55120 42712
rect 55068 42669 55077 42703
rect 55077 42669 55111 42703
rect 55111 42669 55120 42703
rect 55068 42660 55120 42669
rect 12130 42463 12182 42472
rect 12130 42429 12139 42463
rect 12139 42429 12173 42463
rect 12173 42429 12182 42463
rect 12130 42420 12182 42429
rect 55068 42463 55120 42472
rect 55068 42429 55077 42463
rect 55077 42429 55111 42463
rect 55111 42429 55120 42463
rect 55068 42420 55120 42429
rect 12130 41913 12182 41922
rect 12130 41879 12139 41913
rect 12139 41879 12173 41913
rect 12173 41879 12182 41913
rect 12130 41870 12182 41879
rect 55068 41913 55120 41922
rect 55068 41879 55077 41913
rect 55077 41879 55111 41913
rect 55111 41879 55120 41913
rect 55068 41870 55120 41879
rect 12130 41673 12182 41682
rect 12130 41639 12139 41673
rect 12139 41639 12173 41673
rect 12173 41639 12182 41673
rect 12130 41630 12182 41639
rect 55068 41673 55120 41682
rect 55068 41639 55077 41673
rect 55077 41639 55111 41673
rect 55111 41639 55120 41673
rect 55068 41630 55120 41639
rect 12130 41123 12182 41132
rect 12130 41089 12139 41123
rect 12139 41089 12173 41123
rect 12173 41089 12182 41123
rect 12130 41080 12182 41089
rect 55068 41123 55120 41132
rect 55068 41089 55077 41123
rect 55077 41089 55111 41123
rect 55111 41089 55120 41123
rect 55068 41080 55120 41089
rect 12130 40883 12182 40892
rect 12130 40849 12139 40883
rect 12139 40849 12173 40883
rect 12173 40849 12182 40883
rect 12130 40840 12182 40849
rect 55068 40883 55120 40892
rect 55068 40849 55077 40883
rect 55077 40849 55111 40883
rect 55111 40849 55120 40883
rect 55068 40840 55120 40849
rect 12130 40333 12182 40342
rect 12130 40299 12139 40333
rect 12139 40299 12173 40333
rect 12173 40299 12182 40333
rect 12130 40290 12182 40299
rect 55068 40333 55120 40342
rect 55068 40299 55077 40333
rect 55077 40299 55111 40333
rect 55111 40299 55120 40333
rect 55068 40290 55120 40299
rect 12130 40093 12182 40102
rect 12130 40059 12139 40093
rect 12139 40059 12173 40093
rect 12173 40059 12182 40093
rect 12130 40050 12182 40059
rect 55068 40093 55120 40102
rect 55068 40059 55077 40093
rect 55077 40059 55111 40093
rect 55111 40059 55120 40093
rect 55068 40050 55120 40059
rect 12130 39543 12182 39552
rect 12130 39509 12139 39543
rect 12139 39509 12173 39543
rect 12173 39509 12182 39543
rect 12130 39500 12182 39509
rect 55068 39543 55120 39552
rect 55068 39509 55077 39543
rect 55077 39509 55111 39543
rect 55111 39509 55120 39543
rect 55068 39500 55120 39509
rect 12130 39303 12182 39312
rect 12130 39269 12139 39303
rect 12139 39269 12173 39303
rect 12173 39269 12182 39303
rect 12130 39260 12182 39269
rect 55068 39303 55120 39312
rect 55068 39269 55077 39303
rect 55077 39269 55111 39303
rect 55111 39269 55120 39303
rect 55068 39260 55120 39269
rect 12130 38753 12182 38762
rect 12130 38719 12139 38753
rect 12139 38719 12173 38753
rect 12173 38719 12182 38753
rect 12130 38710 12182 38719
rect 55068 38753 55120 38762
rect 55068 38719 55077 38753
rect 55077 38719 55111 38753
rect 55111 38719 55120 38753
rect 55068 38710 55120 38719
rect 12130 38513 12182 38522
rect 12130 38479 12139 38513
rect 12139 38479 12173 38513
rect 12173 38479 12182 38513
rect 12130 38470 12182 38479
rect 55068 38513 55120 38522
rect 55068 38479 55077 38513
rect 55077 38479 55111 38513
rect 55111 38479 55120 38513
rect 55068 38470 55120 38479
rect 12130 37963 12182 37972
rect 12130 37929 12139 37963
rect 12139 37929 12173 37963
rect 12173 37929 12182 37963
rect 12130 37920 12182 37929
rect 55068 37963 55120 37972
rect 55068 37929 55077 37963
rect 55077 37929 55111 37963
rect 55111 37929 55120 37963
rect 55068 37920 55120 37929
rect 12130 37723 12182 37732
rect 12130 37689 12139 37723
rect 12139 37689 12173 37723
rect 12173 37689 12182 37723
rect 12130 37680 12182 37689
rect 55068 37723 55120 37732
rect 55068 37689 55077 37723
rect 55077 37689 55111 37723
rect 55111 37689 55120 37723
rect 55068 37680 55120 37689
rect 12130 37173 12182 37182
rect 12130 37139 12139 37173
rect 12139 37139 12173 37173
rect 12173 37139 12182 37173
rect 12130 37130 12182 37139
rect 55068 37173 55120 37182
rect 55068 37139 55077 37173
rect 55077 37139 55111 37173
rect 55111 37139 55120 37173
rect 55068 37130 55120 37139
rect 12130 36933 12182 36942
rect 12130 36899 12139 36933
rect 12139 36899 12173 36933
rect 12173 36899 12182 36933
rect 12130 36890 12182 36899
rect 55068 36933 55120 36942
rect 55068 36899 55077 36933
rect 55077 36899 55111 36933
rect 55111 36899 55120 36933
rect 55068 36890 55120 36899
rect 12130 36383 12182 36392
rect 12130 36349 12139 36383
rect 12139 36349 12173 36383
rect 12173 36349 12182 36383
rect 12130 36340 12182 36349
rect 55068 36383 55120 36392
rect 55068 36349 55077 36383
rect 55077 36349 55111 36383
rect 55111 36349 55120 36383
rect 55068 36340 55120 36349
rect 12130 36143 12182 36152
rect 12130 36109 12139 36143
rect 12139 36109 12173 36143
rect 12173 36109 12182 36143
rect 12130 36100 12182 36109
rect 55068 36143 55120 36152
rect 55068 36109 55077 36143
rect 55077 36109 55111 36143
rect 55111 36109 55120 36143
rect 55068 36100 55120 36109
rect 12130 35593 12182 35602
rect 12130 35559 12139 35593
rect 12139 35559 12173 35593
rect 12173 35559 12182 35593
rect 12130 35550 12182 35559
rect 55068 35593 55120 35602
rect 55068 35559 55077 35593
rect 55077 35559 55111 35593
rect 55111 35559 55120 35593
rect 55068 35550 55120 35559
rect 12130 35353 12182 35362
rect 12130 35319 12139 35353
rect 12139 35319 12173 35353
rect 12173 35319 12182 35353
rect 12130 35310 12182 35319
rect 55068 35353 55120 35362
rect 55068 35319 55077 35353
rect 55077 35319 55111 35353
rect 55111 35319 55120 35353
rect 55068 35310 55120 35319
rect 12130 34803 12182 34812
rect 12130 34769 12139 34803
rect 12139 34769 12173 34803
rect 12173 34769 12182 34803
rect 12130 34760 12182 34769
rect 55068 34803 55120 34812
rect 55068 34769 55077 34803
rect 55077 34769 55111 34803
rect 55111 34769 55120 34803
rect 55068 34760 55120 34769
rect 12130 34563 12182 34572
rect 12130 34529 12139 34563
rect 12139 34529 12173 34563
rect 12173 34529 12182 34563
rect 12130 34520 12182 34529
rect 55068 34563 55120 34572
rect 55068 34529 55077 34563
rect 55077 34529 55111 34563
rect 55111 34529 55120 34563
rect 55068 34520 55120 34529
rect 12130 34013 12182 34022
rect 12130 33979 12139 34013
rect 12139 33979 12173 34013
rect 12173 33979 12182 34013
rect 12130 33970 12182 33979
rect 55068 34013 55120 34022
rect 55068 33979 55077 34013
rect 55077 33979 55111 34013
rect 55111 33979 55120 34013
rect 55068 33970 55120 33979
rect 12130 33773 12182 33782
rect 12130 33739 12139 33773
rect 12139 33739 12173 33773
rect 12173 33739 12182 33773
rect 12130 33730 12182 33739
rect 55068 33773 55120 33782
rect 55068 33739 55077 33773
rect 55077 33739 55111 33773
rect 55111 33739 55120 33773
rect 55068 33730 55120 33739
rect 12130 33223 12182 33232
rect 12130 33189 12139 33223
rect 12139 33189 12173 33223
rect 12173 33189 12182 33223
rect 12130 33180 12182 33189
rect 55068 33223 55120 33232
rect 55068 33189 55077 33223
rect 55077 33189 55111 33223
rect 55111 33189 55120 33223
rect 55068 33180 55120 33189
rect 12130 32983 12182 32992
rect 12130 32949 12139 32983
rect 12139 32949 12173 32983
rect 12173 32949 12182 32983
rect 12130 32940 12182 32949
rect 55068 32983 55120 32992
rect 55068 32949 55077 32983
rect 55077 32949 55111 32983
rect 55111 32949 55120 32983
rect 55068 32940 55120 32949
rect 12130 32433 12182 32442
rect 12130 32399 12139 32433
rect 12139 32399 12173 32433
rect 12173 32399 12182 32433
rect 12130 32390 12182 32399
rect 55068 32433 55120 32442
rect 55068 32399 55077 32433
rect 55077 32399 55111 32433
rect 55111 32399 55120 32433
rect 55068 32390 55120 32399
rect 12130 32193 12182 32202
rect 12130 32159 12139 32193
rect 12139 32159 12173 32193
rect 12173 32159 12182 32193
rect 12130 32150 12182 32159
rect 55068 32193 55120 32202
rect 55068 32159 55077 32193
rect 55077 32159 55111 32193
rect 55111 32159 55120 32193
rect 55068 32150 55120 32159
rect 12130 31643 12182 31652
rect 12130 31609 12139 31643
rect 12139 31609 12173 31643
rect 12173 31609 12182 31643
rect 12130 31600 12182 31609
rect 55068 31643 55120 31652
rect 55068 31609 55077 31643
rect 55077 31609 55111 31643
rect 55111 31609 55120 31643
rect 55068 31600 55120 31609
rect 12130 31403 12182 31412
rect 12130 31369 12139 31403
rect 12139 31369 12173 31403
rect 12173 31369 12182 31403
rect 12130 31360 12182 31369
rect 55068 31403 55120 31412
rect 55068 31369 55077 31403
rect 55077 31369 55111 31403
rect 55111 31369 55120 31403
rect 55068 31360 55120 31369
rect 12130 30853 12182 30862
rect 12130 30819 12139 30853
rect 12139 30819 12173 30853
rect 12173 30819 12182 30853
rect 12130 30810 12182 30819
rect 55068 30853 55120 30862
rect 55068 30819 55077 30853
rect 55077 30819 55111 30853
rect 55111 30819 55120 30853
rect 55068 30810 55120 30819
rect 12130 30613 12182 30622
rect 12130 30579 12139 30613
rect 12139 30579 12173 30613
rect 12173 30579 12182 30613
rect 12130 30570 12182 30579
rect 55068 30613 55120 30622
rect 55068 30579 55077 30613
rect 55077 30579 55111 30613
rect 55111 30579 55120 30613
rect 55068 30570 55120 30579
rect 12130 30063 12182 30072
rect 12130 30029 12139 30063
rect 12139 30029 12173 30063
rect 12173 30029 12182 30063
rect 12130 30020 12182 30029
rect 55068 30063 55120 30072
rect 55068 30029 55077 30063
rect 55077 30029 55111 30063
rect 55111 30029 55120 30063
rect 55068 30020 55120 30029
rect 12130 29823 12182 29832
rect 12130 29789 12139 29823
rect 12139 29789 12173 29823
rect 12173 29789 12182 29823
rect 12130 29780 12182 29789
rect 55068 29823 55120 29832
rect 55068 29789 55077 29823
rect 55077 29789 55111 29823
rect 55111 29789 55120 29823
rect 55068 29780 55120 29789
rect 12130 29273 12182 29282
rect 12130 29239 12139 29273
rect 12139 29239 12173 29273
rect 12173 29239 12182 29273
rect 12130 29230 12182 29239
rect 55068 29273 55120 29282
rect 55068 29239 55077 29273
rect 55077 29239 55111 29273
rect 55111 29239 55120 29273
rect 55068 29230 55120 29239
rect 12130 29033 12182 29042
rect 12130 28999 12139 29033
rect 12139 28999 12173 29033
rect 12173 28999 12182 29033
rect 12130 28990 12182 28999
rect 55068 29033 55120 29042
rect 55068 28999 55077 29033
rect 55077 28999 55111 29033
rect 55111 28999 55120 29033
rect 55068 28990 55120 28999
rect 12130 28483 12182 28492
rect 12130 28449 12139 28483
rect 12139 28449 12173 28483
rect 12173 28449 12182 28483
rect 12130 28440 12182 28449
rect 55068 28483 55120 28492
rect 55068 28449 55077 28483
rect 55077 28449 55111 28483
rect 55111 28449 55120 28483
rect 55068 28440 55120 28449
rect 12130 28243 12182 28252
rect 12130 28209 12139 28243
rect 12139 28209 12173 28243
rect 12173 28209 12182 28243
rect 12130 28200 12182 28209
rect 55068 28243 55120 28252
rect 55068 28209 55077 28243
rect 55077 28209 55111 28243
rect 55111 28209 55120 28243
rect 55068 28200 55120 28209
rect 12130 27693 12182 27702
rect 12130 27659 12139 27693
rect 12139 27659 12173 27693
rect 12173 27659 12182 27693
rect 12130 27650 12182 27659
rect 55068 27693 55120 27702
rect 55068 27659 55077 27693
rect 55077 27659 55111 27693
rect 55111 27659 55120 27693
rect 55068 27650 55120 27659
rect 12130 27453 12182 27462
rect 12130 27419 12139 27453
rect 12139 27419 12173 27453
rect 12173 27419 12182 27453
rect 12130 27410 12182 27419
rect 55068 27453 55120 27462
rect 55068 27419 55077 27453
rect 55077 27419 55111 27453
rect 55111 27419 55120 27453
rect 55068 27410 55120 27419
rect 12130 26903 12182 26912
rect 12130 26869 12139 26903
rect 12139 26869 12173 26903
rect 12173 26869 12182 26903
rect 12130 26860 12182 26869
rect 55068 26903 55120 26912
rect 55068 26869 55077 26903
rect 55077 26869 55111 26903
rect 55111 26869 55120 26903
rect 55068 26860 55120 26869
rect 12130 26663 12182 26672
rect 12130 26629 12139 26663
rect 12139 26629 12173 26663
rect 12173 26629 12182 26663
rect 12130 26620 12182 26629
rect 55068 26663 55120 26672
rect 55068 26629 55077 26663
rect 55077 26629 55111 26663
rect 55111 26629 55120 26663
rect 55068 26620 55120 26629
rect 12130 26113 12182 26122
rect 12130 26079 12139 26113
rect 12139 26079 12173 26113
rect 12173 26079 12182 26113
rect 12130 26070 12182 26079
rect 55068 26113 55120 26122
rect 55068 26079 55077 26113
rect 55077 26079 55111 26113
rect 55111 26079 55120 26113
rect 55068 26070 55120 26079
rect 12130 25873 12182 25882
rect 12130 25839 12139 25873
rect 12139 25839 12173 25873
rect 12173 25839 12182 25873
rect 12130 25830 12182 25839
rect 55068 25873 55120 25882
rect 55068 25839 55077 25873
rect 55077 25839 55111 25873
rect 55111 25839 55120 25873
rect 55068 25830 55120 25839
rect 12130 25323 12182 25332
rect 12130 25289 12139 25323
rect 12139 25289 12173 25323
rect 12173 25289 12182 25323
rect 12130 25280 12182 25289
rect 55068 25323 55120 25332
rect 55068 25289 55077 25323
rect 55077 25289 55111 25323
rect 55111 25289 55120 25323
rect 55068 25280 55120 25289
rect 12130 25083 12182 25092
rect 12130 25049 12139 25083
rect 12139 25049 12173 25083
rect 12173 25049 12182 25083
rect 12130 25040 12182 25049
rect 55068 25083 55120 25092
rect 55068 25049 55077 25083
rect 55077 25049 55111 25083
rect 55111 25049 55120 25083
rect 55068 25040 55120 25049
rect 12130 24533 12182 24542
rect 12130 24499 12139 24533
rect 12139 24499 12173 24533
rect 12173 24499 12182 24533
rect 12130 24490 12182 24499
rect 55068 24533 55120 24542
rect 55068 24499 55077 24533
rect 55077 24499 55111 24533
rect 55111 24499 55120 24533
rect 55068 24490 55120 24499
rect 12130 24293 12182 24302
rect 12130 24259 12139 24293
rect 12139 24259 12173 24293
rect 12173 24259 12182 24293
rect 12130 24250 12182 24259
rect 55068 24293 55120 24302
rect 55068 24259 55077 24293
rect 55077 24259 55111 24293
rect 55111 24259 55120 24293
rect 55068 24250 55120 24259
rect 12130 23743 12182 23752
rect 12130 23709 12139 23743
rect 12139 23709 12173 23743
rect 12173 23709 12182 23743
rect 12130 23700 12182 23709
rect 55068 23743 55120 23752
rect 55068 23709 55077 23743
rect 55077 23709 55111 23743
rect 55111 23709 55120 23743
rect 55068 23700 55120 23709
rect 12130 23503 12182 23512
rect 12130 23469 12139 23503
rect 12139 23469 12173 23503
rect 12173 23469 12182 23503
rect 12130 23460 12182 23469
rect 55068 23503 55120 23512
rect 55068 23469 55077 23503
rect 55077 23469 55111 23503
rect 55111 23469 55120 23503
rect 55068 23460 55120 23469
rect 12130 22953 12182 22962
rect 12130 22919 12139 22953
rect 12139 22919 12173 22953
rect 12173 22919 12182 22953
rect 12130 22910 12182 22919
rect 55068 22953 55120 22962
rect 55068 22919 55077 22953
rect 55077 22919 55111 22953
rect 55111 22919 55120 22953
rect 55068 22910 55120 22919
rect 12130 22713 12182 22722
rect 12130 22679 12139 22713
rect 12139 22679 12173 22713
rect 12173 22679 12182 22713
rect 12130 22670 12182 22679
rect 55068 22713 55120 22722
rect 55068 22679 55077 22713
rect 55077 22679 55111 22713
rect 55111 22679 55120 22713
rect 55068 22670 55120 22679
rect 12130 22163 12182 22172
rect 12130 22129 12139 22163
rect 12139 22129 12173 22163
rect 12173 22129 12182 22163
rect 12130 22120 12182 22129
rect 55068 22163 55120 22172
rect 55068 22129 55077 22163
rect 55077 22129 55111 22163
rect 55111 22129 55120 22163
rect 55068 22120 55120 22129
rect 12130 21923 12182 21932
rect 12130 21889 12139 21923
rect 12139 21889 12173 21923
rect 12173 21889 12182 21923
rect 12130 21880 12182 21889
rect 55068 21923 55120 21932
rect 55068 21889 55077 21923
rect 55077 21889 55111 21923
rect 55111 21889 55120 21923
rect 55068 21880 55120 21889
rect 12130 21373 12182 21382
rect 12130 21339 12139 21373
rect 12139 21339 12173 21373
rect 12173 21339 12182 21373
rect 12130 21330 12182 21339
rect 55068 21373 55120 21382
rect 55068 21339 55077 21373
rect 55077 21339 55111 21373
rect 55111 21339 55120 21373
rect 55068 21330 55120 21339
rect 12130 21133 12182 21142
rect 12130 21099 12139 21133
rect 12139 21099 12173 21133
rect 12173 21099 12182 21133
rect 12130 21090 12182 21099
rect 55068 21133 55120 21142
rect 55068 21099 55077 21133
rect 55077 21099 55111 21133
rect 55111 21099 55120 21133
rect 55068 21090 55120 21099
rect 12130 20583 12182 20592
rect 12130 20549 12139 20583
rect 12139 20549 12173 20583
rect 12173 20549 12182 20583
rect 12130 20540 12182 20549
rect 55068 20583 55120 20592
rect 55068 20549 55077 20583
rect 55077 20549 55111 20583
rect 55111 20549 55120 20583
rect 55068 20540 55120 20549
rect 12130 20343 12182 20352
rect 12130 20309 12139 20343
rect 12139 20309 12173 20343
rect 12173 20309 12182 20343
rect 12130 20300 12182 20309
rect 55068 20343 55120 20352
rect 55068 20309 55077 20343
rect 55077 20309 55111 20343
rect 55111 20309 55120 20343
rect 55068 20300 55120 20309
rect 12130 19793 12182 19802
rect 12130 19759 12139 19793
rect 12139 19759 12173 19793
rect 12173 19759 12182 19793
rect 12130 19750 12182 19759
rect 55068 19793 55120 19802
rect 55068 19759 55077 19793
rect 55077 19759 55111 19793
rect 55111 19759 55120 19793
rect 55068 19750 55120 19759
rect 12130 19553 12182 19562
rect 12130 19519 12139 19553
rect 12139 19519 12173 19553
rect 12173 19519 12182 19553
rect 12130 19510 12182 19519
rect 55068 19553 55120 19562
rect 55068 19519 55077 19553
rect 55077 19519 55111 19553
rect 55111 19519 55120 19553
rect 55068 19510 55120 19519
rect 12130 19003 12182 19012
rect 12130 18969 12139 19003
rect 12139 18969 12173 19003
rect 12173 18969 12182 19003
rect 12130 18960 12182 18969
rect 55068 19003 55120 19012
rect 55068 18969 55077 19003
rect 55077 18969 55111 19003
rect 55111 18969 55120 19003
rect 55068 18960 55120 18969
rect 12130 18763 12182 18772
rect 12130 18729 12139 18763
rect 12139 18729 12173 18763
rect 12173 18729 12182 18763
rect 12130 18720 12182 18729
rect 55068 18763 55120 18772
rect 55068 18729 55077 18763
rect 55077 18729 55111 18763
rect 55111 18729 55120 18763
rect 55068 18720 55120 18729
rect 12130 18213 12182 18222
rect 12130 18179 12139 18213
rect 12139 18179 12173 18213
rect 12173 18179 12182 18213
rect 12130 18170 12182 18179
rect 55068 18213 55120 18222
rect 55068 18179 55077 18213
rect 55077 18179 55111 18213
rect 55111 18179 55120 18213
rect 55068 18170 55120 18179
rect 12130 17973 12182 17982
rect 12130 17939 12139 17973
rect 12139 17939 12173 17973
rect 12173 17939 12182 17973
rect 12130 17930 12182 17939
rect 55068 17973 55120 17982
rect 55068 17939 55077 17973
rect 55077 17939 55111 17973
rect 55111 17939 55120 17973
rect 55068 17930 55120 17939
rect 12130 17423 12182 17432
rect 12130 17389 12139 17423
rect 12139 17389 12173 17423
rect 12173 17389 12182 17423
rect 12130 17380 12182 17389
rect 55068 17423 55120 17432
rect 55068 17389 55077 17423
rect 55077 17389 55111 17423
rect 55111 17389 55120 17423
rect 55068 17380 55120 17389
rect 12130 17183 12182 17192
rect 12130 17149 12139 17183
rect 12139 17149 12173 17183
rect 12173 17149 12182 17183
rect 12130 17140 12182 17149
rect 55068 17183 55120 17192
rect 55068 17149 55077 17183
rect 55077 17149 55111 17183
rect 55111 17149 55120 17183
rect 55068 17140 55120 17149
rect 12130 16633 12182 16642
rect 12130 16599 12139 16633
rect 12139 16599 12173 16633
rect 12173 16599 12182 16633
rect 12130 16590 12182 16599
rect 55068 16633 55120 16642
rect 55068 16599 55077 16633
rect 55077 16599 55111 16633
rect 55111 16599 55120 16633
rect 55068 16590 55120 16599
rect 12130 16393 12182 16402
rect 12130 16359 12139 16393
rect 12139 16359 12173 16393
rect 12173 16359 12182 16393
rect 12130 16350 12182 16359
rect 55068 16393 55120 16402
rect 55068 16359 55077 16393
rect 55077 16359 55111 16393
rect 55111 16359 55120 16393
rect 55068 16350 55120 16359
rect 12130 15843 12182 15852
rect 12130 15809 12139 15843
rect 12139 15809 12173 15843
rect 12173 15809 12182 15843
rect 12130 15800 12182 15809
rect 55068 15843 55120 15852
rect 55068 15809 55077 15843
rect 55077 15809 55111 15843
rect 55111 15809 55120 15843
rect 55068 15800 55120 15809
rect 12130 15603 12182 15612
rect 12130 15569 12139 15603
rect 12139 15569 12173 15603
rect 12173 15569 12182 15603
rect 12130 15560 12182 15569
rect 55068 15603 55120 15612
rect 55068 15569 55077 15603
rect 55077 15569 55111 15603
rect 55111 15569 55120 15603
rect 55068 15560 55120 15569
rect 12130 15053 12182 15062
rect 12130 15019 12139 15053
rect 12139 15019 12173 15053
rect 12173 15019 12182 15053
rect 12130 15010 12182 15019
rect 55068 15053 55120 15062
rect 55068 15019 55077 15053
rect 55077 15019 55111 15053
rect 55111 15019 55120 15053
rect 55068 15010 55120 15019
rect 12130 14813 12182 14822
rect 12130 14779 12139 14813
rect 12139 14779 12173 14813
rect 12173 14779 12182 14813
rect 12130 14770 12182 14779
rect 55068 14813 55120 14822
rect 55068 14779 55077 14813
rect 55077 14779 55111 14813
rect 55111 14779 55120 14813
rect 55068 14770 55120 14779
rect 12130 14263 12182 14272
rect 12130 14229 12139 14263
rect 12139 14229 12173 14263
rect 12173 14229 12182 14263
rect 12130 14220 12182 14229
rect 55068 14263 55120 14272
rect 55068 14229 55077 14263
rect 55077 14229 55111 14263
rect 55111 14229 55120 14263
rect 55068 14220 55120 14229
rect 12130 14023 12182 14032
rect 12130 13989 12139 14023
rect 12139 13989 12173 14023
rect 12173 13989 12182 14023
rect 12130 13980 12182 13989
rect 55068 14023 55120 14032
rect 55068 13989 55077 14023
rect 55077 13989 55111 14023
rect 55111 13989 55120 14023
rect 55068 13980 55120 13989
rect 12130 13473 12182 13482
rect 12130 13439 12139 13473
rect 12139 13439 12173 13473
rect 12173 13439 12182 13473
rect 12130 13430 12182 13439
rect 55068 13473 55120 13482
rect 55068 13439 55077 13473
rect 55077 13439 55111 13473
rect 55111 13439 55120 13473
rect 55068 13430 55120 13439
rect 12130 13233 12182 13242
rect 12130 13199 12139 13233
rect 12139 13199 12173 13233
rect 12173 13199 12182 13233
rect 12130 13190 12182 13199
rect 55068 13233 55120 13242
rect 55068 13199 55077 13233
rect 55077 13199 55111 13233
rect 55111 13199 55120 13233
rect 55068 13190 55120 13199
rect 12130 12683 12182 12692
rect 12130 12649 12139 12683
rect 12139 12649 12173 12683
rect 12173 12649 12182 12683
rect 12130 12640 12182 12649
rect 55068 12683 55120 12692
rect 55068 12649 55077 12683
rect 55077 12649 55111 12683
rect 55111 12649 55120 12683
rect 55068 12640 55120 12649
rect 12130 12443 12182 12452
rect 12130 12409 12139 12443
rect 12139 12409 12173 12443
rect 12173 12409 12182 12443
rect 12130 12400 12182 12409
rect 55068 12443 55120 12452
rect 55068 12409 55077 12443
rect 55077 12409 55111 12443
rect 55111 12409 55120 12443
rect 55068 12400 55120 12409
rect 12130 11893 12182 11902
rect 12130 11859 12139 11893
rect 12139 11859 12173 11893
rect 12173 11859 12182 11893
rect 12130 11850 12182 11859
rect 55068 11893 55120 11902
rect 55068 11859 55077 11893
rect 55077 11859 55111 11893
rect 55111 11859 55120 11893
rect 55068 11850 55120 11859
rect 12130 11653 12182 11662
rect 12130 11619 12139 11653
rect 12139 11619 12173 11653
rect 12173 11619 12182 11653
rect 12130 11610 12182 11619
rect 55068 11653 55120 11662
rect 55068 11619 55077 11653
rect 55077 11619 55111 11653
rect 55111 11619 55120 11653
rect 55068 11610 55120 11619
rect 12130 11103 12182 11112
rect 12130 11069 12139 11103
rect 12139 11069 12173 11103
rect 12173 11069 12182 11103
rect 12130 11060 12182 11069
rect 55068 11103 55120 11112
rect 55068 11069 55077 11103
rect 55077 11069 55111 11103
rect 55111 11069 55120 11103
rect 55068 11060 55120 11069
rect 12130 10863 12182 10872
rect 12130 10829 12139 10863
rect 12139 10829 12173 10863
rect 12173 10829 12182 10863
rect 12130 10820 12182 10829
rect 55068 10863 55120 10872
rect 55068 10829 55077 10863
rect 55077 10829 55111 10863
rect 55111 10829 55120 10863
rect 55068 10820 55120 10829
rect 12130 10313 12182 10322
rect 12130 10279 12139 10313
rect 12139 10279 12173 10313
rect 12173 10279 12182 10313
rect 12130 10270 12182 10279
rect 55068 10313 55120 10322
rect 55068 10279 55077 10313
rect 55077 10279 55111 10313
rect 55111 10279 55120 10313
rect 55068 10270 55120 10279
rect 12130 10073 12182 10082
rect 12130 10039 12139 10073
rect 12139 10039 12173 10073
rect 12173 10039 12182 10073
rect 12130 10030 12182 10039
rect 13551 8230 13603 8282
rect 6731 7652 6783 7661
rect 6731 7618 6740 7652
rect 6740 7618 6774 7652
rect 6774 7618 6783 7652
rect 6731 7609 6783 7618
rect 7130 6945 7182 6954
rect 7130 6911 7139 6945
rect 7139 6911 7173 6945
rect 7173 6911 7182 6945
rect 7130 6902 7182 6911
rect 6731 6238 6783 6247
rect 6731 6204 6740 6238
rect 6740 6204 6774 6238
rect 6774 6204 6783 6238
rect 6731 6195 6783 6204
rect 7130 5531 7182 5540
rect 7130 5497 7139 5531
rect 7139 5497 7173 5531
rect 7173 5497 7182 5531
rect 7130 5488 7182 5497
rect 6731 4824 6783 4833
rect 6731 4790 6740 4824
rect 6740 4790 6774 4824
rect 6774 4790 6783 4824
rect 6731 4781 6783 4790
<< metal2 >>
rect 55277 65071 55305 67312
rect 55263 65062 55319 65071
rect 55263 64997 55319 65006
rect 53645 62684 53701 62693
rect 53645 62619 53701 62628
rect 55277 61526 55305 64997
rect 55401 62544 55429 67312
rect 60341 66133 60397 66142
rect 60341 66068 60397 66077
rect 59337 65426 59393 65435
rect 59337 65361 59393 65370
rect 59942 65426 59998 65435
rect 59942 65361 59998 65370
rect 59351 64355 59379 65361
rect 60341 64719 60397 64728
rect 60341 64654 60397 64663
rect 59337 64346 59393 64355
rect 59337 64281 59393 64290
rect 59201 64222 59257 64231
rect 59201 64157 59257 64166
rect 59215 64021 59243 64157
rect 59201 64012 59257 64021
rect 59201 63947 59257 63956
rect 59942 64012 59998 64021
rect 59942 63947 59998 63956
rect 60341 63305 60397 63314
rect 60341 63240 60397 63249
rect 55387 62535 55443 62544
rect 55387 62470 55443 62479
rect 55401 61526 55429 62470
rect 59262 61021 59290 61049
rect 55068 60882 55120 60888
rect 54967 60849 55068 60877
rect 55068 60824 55120 60830
rect 12130 60642 12182 60648
rect 55068 60642 55120 60648
rect 54967 60595 55068 60623
rect 12130 60584 12182 60590
rect 55068 60584 55120 60590
rect 12142 60403 12170 60584
rect 12142 60375 12283 60403
rect 12142 60279 12283 60307
rect 12142 60098 12170 60279
rect 12130 60092 12182 60098
rect 55068 60092 55120 60098
rect 54967 60059 55068 60087
rect 12130 60034 12182 60040
rect 55068 60034 55120 60040
rect 12130 59852 12182 59858
rect 55068 59852 55120 59858
rect 54967 59805 55068 59833
rect 12130 59794 12182 59800
rect 55068 59794 55120 59800
rect 12142 59613 12170 59794
rect 12142 59585 12283 59613
rect 12142 59489 12283 59517
rect 12142 59308 12170 59489
rect 12130 59302 12182 59308
rect 55068 59302 55120 59308
rect 54967 59269 55068 59297
rect 12130 59244 12182 59250
rect 55068 59244 55120 59250
rect 12130 59062 12182 59068
rect 55068 59062 55120 59068
rect 54967 59015 55068 59043
rect 12130 59004 12182 59010
rect 55068 59004 55120 59010
rect 12142 58823 12170 59004
rect 12142 58795 12283 58823
rect 12142 58699 12283 58727
rect 12142 58518 12170 58699
rect 12130 58512 12182 58518
rect 55068 58512 55120 58518
rect 54967 58479 55068 58507
rect 12130 58454 12182 58460
rect 55068 58454 55120 58460
rect 12130 58272 12182 58278
rect 55068 58272 55120 58278
rect 54967 58225 55068 58253
rect 12130 58214 12182 58220
rect 55068 58214 55120 58220
rect 12142 58033 12170 58214
rect 12142 58005 12283 58033
rect 12142 57909 12283 57937
rect 12142 57728 12170 57909
rect 12130 57722 12182 57728
rect 55068 57722 55120 57728
rect 54967 57689 55068 57717
rect 12130 57664 12182 57670
rect 55068 57664 55120 57670
rect 12130 57482 12182 57488
rect 55068 57482 55120 57488
rect 54967 57435 55068 57463
rect 12130 57424 12182 57430
rect 55068 57424 55120 57430
rect 12142 57243 12170 57424
rect 12142 57215 12283 57243
rect 12142 57119 12283 57147
rect 12142 56938 12170 57119
rect 12130 56932 12182 56938
rect 55068 56932 55120 56938
rect 54967 56899 55068 56927
rect 12130 56874 12182 56880
rect 55068 56874 55120 56880
rect 12130 56692 12182 56698
rect 55068 56692 55120 56698
rect 54967 56645 55068 56673
rect 12130 56634 12182 56640
rect 55068 56634 55120 56640
rect 12142 56453 12170 56634
rect 12142 56425 12283 56453
rect 12142 56329 12283 56357
rect 12142 56148 12170 56329
rect 12130 56142 12182 56148
rect 55068 56142 55120 56148
rect 54967 56109 55068 56137
rect 12130 56084 12182 56090
rect 55068 56084 55120 56090
rect 12130 55902 12182 55908
rect 55068 55902 55120 55908
rect 54967 55855 55068 55883
rect 12130 55844 12182 55850
rect 55068 55844 55120 55850
rect 12142 55663 12170 55844
rect 12142 55635 12283 55663
rect 12142 55539 12283 55567
rect 12142 55358 12170 55539
rect 12130 55352 12182 55358
rect 55068 55352 55120 55358
rect 54967 55319 55068 55347
rect 12130 55294 12182 55300
rect 55068 55294 55120 55300
rect 12130 55112 12182 55118
rect 55068 55112 55120 55118
rect 54967 55065 55068 55093
rect 12130 55054 12182 55060
rect 55068 55054 55120 55060
rect 12142 54873 12170 55054
rect 12142 54845 12283 54873
rect 12142 54749 12283 54777
rect 12142 54568 12170 54749
rect 12130 54562 12182 54568
rect 55068 54562 55120 54568
rect 54967 54529 55068 54557
rect 12130 54504 12182 54510
rect 55068 54504 55120 54510
rect 12130 54322 12182 54328
rect 55068 54322 55120 54328
rect 54967 54275 55068 54303
rect 12130 54264 12182 54270
rect 55068 54264 55120 54270
rect 12142 54083 12170 54264
rect 12142 54055 12283 54083
rect 12142 53959 12283 53987
rect 12142 53778 12170 53959
rect 12130 53772 12182 53778
rect 55068 53772 55120 53778
rect 54967 53739 55068 53767
rect 12130 53714 12182 53720
rect 55068 53714 55120 53720
rect 12130 53532 12182 53538
rect 55068 53532 55120 53538
rect 54967 53485 55068 53513
rect 12130 53474 12182 53480
rect 55068 53474 55120 53480
rect 12142 53293 12170 53474
rect 12142 53265 12283 53293
rect 12142 53169 12283 53197
rect 12142 52988 12170 53169
rect 12130 52982 12182 52988
rect 55068 52982 55120 52988
rect 54967 52949 55068 52977
rect 12130 52924 12182 52930
rect 55068 52924 55120 52930
rect 12130 52742 12182 52748
rect 55068 52742 55120 52748
rect 54967 52695 55068 52723
rect 12130 52684 12182 52690
rect 55068 52684 55120 52690
rect 12142 52503 12170 52684
rect 12142 52475 12283 52503
rect 12142 52379 12283 52407
rect 12142 52198 12170 52379
rect 12130 52192 12182 52198
rect 55068 52192 55120 52198
rect 54967 52159 55068 52187
rect 12130 52134 12182 52140
rect 55068 52134 55120 52140
rect 12130 51952 12182 51958
rect 55068 51952 55120 51958
rect 54967 51905 55068 51933
rect 12130 51894 12182 51900
rect 55068 51894 55120 51900
rect 12142 51713 12170 51894
rect 12142 51685 12283 51713
rect 12142 51589 12283 51617
rect 12142 51408 12170 51589
rect 12130 51402 12182 51408
rect 55068 51402 55120 51408
rect 54967 51369 55068 51397
rect 12130 51344 12182 51350
rect 55068 51344 55120 51350
rect 12130 51162 12182 51168
rect 55068 51162 55120 51168
rect 54967 51115 55068 51143
rect 12130 51104 12182 51110
rect 55068 51104 55120 51110
rect 12142 50923 12170 51104
rect 12142 50895 12283 50923
rect 12142 50799 12283 50827
rect 12142 50618 12170 50799
rect 12130 50612 12182 50618
rect 55068 50612 55120 50618
rect 54967 50579 55068 50607
rect 12130 50554 12182 50560
rect 55068 50554 55120 50560
rect 12130 50372 12182 50378
rect 55068 50372 55120 50378
rect 54967 50325 55068 50353
rect 12130 50314 12182 50320
rect 55068 50314 55120 50320
rect 12142 50133 12170 50314
rect 12142 50105 12283 50133
rect 12142 50009 12283 50037
rect 12142 49828 12170 50009
rect 12130 49822 12182 49828
rect 55068 49822 55120 49828
rect 54967 49789 55068 49817
rect 12130 49764 12182 49770
rect 55068 49764 55120 49770
rect 12130 49582 12182 49588
rect 55068 49582 55120 49588
rect 54967 49535 55068 49563
rect 12130 49524 12182 49530
rect 55068 49524 55120 49530
rect 12142 49343 12170 49524
rect 12142 49315 12283 49343
rect 12142 49219 12283 49247
rect 12142 49038 12170 49219
rect 12130 49032 12182 49038
rect 55068 49032 55120 49038
rect 54967 48999 55068 49027
rect 12130 48974 12182 48980
rect 55068 48974 55120 48980
rect 12130 48792 12182 48798
rect 55068 48792 55120 48798
rect 54967 48745 55068 48773
rect 12130 48734 12182 48740
rect 55068 48734 55120 48740
rect 12142 48553 12170 48734
rect 12142 48525 12283 48553
rect 12142 48429 12283 48457
rect 12142 48248 12170 48429
rect 12130 48242 12182 48248
rect 55068 48242 55120 48248
rect 54967 48209 55068 48237
rect 12130 48184 12182 48190
rect 55068 48184 55120 48190
rect 12130 48002 12182 48008
rect 55068 48002 55120 48008
rect 54967 47955 55068 47983
rect 12130 47944 12182 47950
rect 55068 47944 55120 47950
rect 12142 47763 12170 47944
rect 12142 47735 12283 47763
rect 12142 47639 12283 47667
rect 12142 47458 12170 47639
rect 12130 47452 12182 47458
rect 55068 47452 55120 47458
rect 54967 47419 55068 47447
rect 12130 47394 12182 47400
rect 55068 47394 55120 47400
rect 12130 47212 12182 47218
rect 55068 47212 55120 47218
rect 54967 47165 55068 47193
rect 12130 47154 12182 47160
rect 55068 47154 55120 47160
rect 12142 46973 12170 47154
rect 12142 46945 12283 46973
rect 12142 46849 12283 46877
rect 12142 46668 12170 46849
rect 12130 46662 12182 46668
rect 55068 46662 55120 46668
rect 54967 46629 55068 46657
rect 12130 46604 12182 46610
rect 55068 46604 55120 46610
rect 12130 46422 12182 46428
rect 55068 46422 55120 46428
rect 54967 46375 55068 46403
rect 12130 46364 12182 46370
rect 55068 46364 55120 46370
rect 12142 46183 12170 46364
rect 12142 46155 12283 46183
rect 12142 46059 12283 46087
rect 12142 45878 12170 46059
rect 12130 45872 12182 45878
rect 55068 45872 55120 45878
rect 54967 45839 55068 45867
rect 12130 45814 12182 45820
rect 55068 45814 55120 45820
rect 12130 45632 12182 45638
rect 55068 45632 55120 45638
rect 54967 45585 55068 45613
rect 12130 45574 12182 45580
rect 55068 45574 55120 45580
rect 12142 45393 12170 45574
rect 12142 45365 12283 45393
rect 12142 45269 12283 45297
rect 12142 45088 12170 45269
rect 12130 45082 12182 45088
rect 55068 45082 55120 45088
rect 54967 45049 55068 45077
rect 12130 45024 12182 45030
rect 55068 45024 55120 45030
rect 12130 44842 12182 44848
rect 55068 44842 55120 44848
rect 54967 44795 55068 44823
rect 12130 44784 12182 44790
rect 55068 44784 55120 44790
rect 12142 44603 12170 44784
rect 12142 44575 12283 44603
rect 12142 44479 12283 44507
rect 12142 44298 12170 44479
rect 12130 44292 12182 44298
rect 55068 44292 55120 44298
rect 54967 44259 55068 44287
rect 12130 44234 12182 44240
rect 55068 44234 55120 44240
rect 12130 44052 12182 44058
rect 55068 44052 55120 44058
rect 54967 44005 55068 44033
rect 12130 43994 12182 44000
rect 55068 43994 55120 44000
rect 12142 43813 12170 43994
rect 12142 43785 12283 43813
rect 12142 43689 12283 43717
rect 12142 43508 12170 43689
rect 12130 43502 12182 43508
rect 55068 43502 55120 43508
rect 54967 43469 55068 43497
rect 12130 43444 12182 43450
rect 55068 43444 55120 43450
rect 12130 43262 12182 43268
rect 55068 43262 55120 43268
rect 54967 43215 55068 43243
rect 12130 43204 12182 43210
rect 55068 43204 55120 43210
rect 12142 43023 12170 43204
rect 12142 42995 12283 43023
rect 12142 42899 12283 42927
rect 12142 42718 12170 42899
rect 12130 42712 12182 42718
rect 55068 42712 55120 42718
rect 54967 42679 55068 42707
rect 12130 42654 12182 42660
rect 55068 42654 55120 42660
rect 12130 42472 12182 42478
rect 55068 42472 55120 42478
rect 54967 42425 55068 42453
rect 12130 42414 12182 42420
rect 55068 42414 55120 42420
rect 12142 42233 12170 42414
rect 12142 42205 12283 42233
rect 12142 42109 12283 42137
rect 12142 41928 12170 42109
rect 12130 41922 12182 41928
rect 55068 41922 55120 41928
rect 54967 41889 55068 41917
rect 12130 41864 12182 41870
rect 55068 41864 55120 41870
rect 12130 41682 12182 41688
rect 55068 41682 55120 41688
rect 54967 41635 55068 41663
rect 12130 41624 12182 41630
rect 55068 41624 55120 41630
rect 12142 41443 12170 41624
rect 12142 41415 12283 41443
rect 12142 41319 12283 41347
rect 12142 41138 12170 41319
rect 12130 41132 12182 41138
rect 55068 41132 55120 41138
rect 54967 41099 55068 41127
rect 12130 41074 12182 41080
rect 55068 41074 55120 41080
rect 12130 40892 12182 40898
rect 55068 40892 55120 40898
rect 54967 40845 55068 40873
rect 12130 40834 12182 40840
rect 55068 40834 55120 40840
rect 12142 40653 12170 40834
rect 12142 40625 12283 40653
rect 12142 40529 12283 40557
rect 12142 40348 12170 40529
rect 12130 40342 12182 40348
rect 55068 40342 55120 40348
rect 54967 40309 55068 40337
rect 12130 40284 12182 40290
rect 55068 40284 55120 40290
rect 12130 40102 12182 40108
rect 55068 40102 55120 40108
rect 54967 40055 55068 40083
rect 12130 40044 12182 40050
rect 55068 40044 55120 40050
rect 12142 39863 12170 40044
rect 12142 39835 12283 39863
rect 12142 39739 12283 39767
rect 12142 39558 12170 39739
rect 12130 39552 12182 39558
rect 55068 39552 55120 39558
rect 54967 39519 55068 39547
rect 12130 39494 12182 39500
rect 55068 39494 55120 39500
rect 12130 39312 12182 39318
rect 55068 39312 55120 39318
rect 54967 39265 55068 39293
rect 12130 39254 12182 39260
rect 55068 39254 55120 39260
rect 12142 39073 12170 39254
rect 12142 39045 12283 39073
rect 12142 38949 12283 38977
rect 12142 38768 12170 38949
rect 12130 38762 12182 38768
rect 55068 38762 55120 38768
rect 54967 38729 55068 38757
rect 12130 38704 12182 38710
rect 55068 38704 55120 38710
rect 12130 38522 12182 38528
rect 55068 38522 55120 38528
rect 54967 38475 55068 38503
rect 12130 38464 12182 38470
rect 55068 38464 55120 38470
rect 12142 38283 12170 38464
rect 12142 38255 12283 38283
rect 12142 38159 12283 38187
rect 12142 37978 12170 38159
rect 12130 37972 12182 37978
rect 55068 37972 55120 37978
rect 54967 37939 55068 37967
rect 12130 37914 12182 37920
rect 55068 37914 55120 37920
rect 12130 37732 12182 37738
rect 55068 37732 55120 37738
rect 54967 37685 55068 37713
rect 12130 37674 12182 37680
rect 55068 37674 55120 37680
rect 12142 37493 12170 37674
rect 12142 37465 12283 37493
rect 12142 37369 12283 37397
rect 12142 37188 12170 37369
rect 12130 37182 12182 37188
rect 55068 37182 55120 37188
rect 54967 37149 55068 37177
rect 12130 37124 12182 37130
rect 55068 37124 55120 37130
rect 12130 36942 12182 36948
rect 55068 36942 55120 36948
rect 54967 36895 55068 36923
rect 12130 36884 12182 36890
rect 55068 36884 55120 36890
rect 12142 36703 12170 36884
rect 12142 36675 12283 36703
rect 12142 36579 12283 36607
rect 12142 36398 12170 36579
rect 12130 36392 12182 36398
rect 55068 36392 55120 36398
rect 54967 36359 55068 36387
rect 12130 36334 12182 36340
rect 55068 36334 55120 36340
rect 12130 36152 12182 36158
rect 55068 36152 55120 36158
rect 54967 36105 55068 36133
rect 12130 36094 12182 36100
rect 55068 36094 55120 36100
rect 12142 35913 12170 36094
rect 12142 35885 12283 35913
rect 12142 35789 12283 35817
rect 12142 35608 12170 35789
rect 12130 35602 12182 35608
rect 55068 35602 55120 35608
rect 54967 35569 55068 35597
rect 12130 35544 12182 35550
rect 55068 35544 55120 35550
rect 12130 35362 12182 35368
rect 55068 35362 55120 35368
rect 54967 35315 55068 35343
rect 12130 35304 12182 35310
rect 55068 35304 55120 35310
rect 12142 35123 12170 35304
rect 12142 35095 12283 35123
rect 12142 34999 12283 35027
rect 12142 34818 12170 34999
rect 12130 34812 12182 34818
rect 55068 34812 55120 34818
rect 54967 34779 55068 34807
rect 12130 34754 12182 34760
rect 55068 34754 55120 34760
rect 12130 34572 12182 34578
rect 55068 34572 55120 34578
rect 54967 34525 55068 34553
rect 12130 34514 12182 34520
rect 55068 34514 55120 34520
rect 12142 34333 12170 34514
rect 12142 34305 12283 34333
rect 12142 34209 12283 34237
rect 12142 34028 12170 34209
rect 12130 34022 12182 34028
rect 55068 34022 55120 34028
rect 54967 33989 55068 34017
rect 12130 33964 12182 33970
rect 55068 33964 55120 33970
rect 12130 33782 12182 33788
rect 55068 33782 55120 33788
rect 54967 33735 55068 33763
rect 12130 33724 12182 33730
rect 55068 33724 55120 33730
rect 12142 33543 12170 33724
rect 12142 33515 12283 33543
rect 12142 33419 12283 33447
rect 12142 33238 12170 33419
rect 12130 33232 12182 33238
rect 55068 33232 55120 33238
rect 54967 33199 55068 33227
rect 12130 33174 12182 33180
rect 55068 33174 55120 33180
rect 12130 32992 12182 32998
rect 55068 32992 55120 32998
rect 54967 32945 55068 32973
rect 12130 32934 12182 32940
rect 55068 32934 55120 32940
rect 12142 32753 12170 32934
rect 12142 32725 12283 32753
rect 12142 32629 12283 32657
rect 12142 32448 12170 32629
rect 12130 32442 12182 32448
rect 55068 32442 55120 32448
rect 54967 32409 55068 32437
rect 12130 32384 12182 32390
rect 55068 32384 55120 32390
rect 12130 32202 12182 32208
rect 55068 32202 55120 32208
rect 54967 32155 55068 32183
rect 12130 32144 12182 32150
rect 55068 32144 55120 32150
rect 12142 31963 12170 32144
rect 12142 31935 12283 31963
rect 12142 31839 12283 31867
rect 12142 31658 12170 31839
rect 12130 31652 12182 31658
rect 55068 31652 55120 31658
rect 54967 31619 55068 31647
rect 12130 31594 12182 31600
rect 55068 31594 55120 31600
rect 12130 31412 12182 31418
rect 55068 31412 55120 31418
rect 54967 31365 55068 31393
rect 12130 31354 12182 31360
rect 55068 31354 55120 31360
rect 12142 31173 12170 31354
rect 12142 31145 12283 31173
rect 12142 31049 12283 31077
rect 12142 30868 12170 31049
rect 12130 30862 12182 30868
rect 55068 30862 55120 30868
rect 54967 30829 55068 30857
rect 12130 30804 12182 30810
rect 55068 30804 55120 30810
rect 12130 30622 12182 30628
rect 55068 30622 55120 30628
rect 54967 30575 55068 30603
rect 12130 30564 12182 30570
rect 55068 30564 55120 30570
rect 12142 30383 12170 30564
rect 12142 30355 12283 30383
rect 12142 30259 12283 30287
rect 12142 30078 12170 30259
rect 12130 30072 12182 30078
rect 55068 30072 55120 30078
rect 54967 30039 55068 30067
rect 12130 30014 12182 30020
rect 55068 30014 55120 30020
rect 12130 29832 12182 29838
rect 55068 29832 55120 29838
rect 54967 29785 55068 29813
rect 12130 29774 12182 29780
rect 55068 29774 55120 29780
rect 12142 29593 12170 29774
rect 12142 29565 12283 29593
rect 12142 29469 12283 29497
rect 12142 29288 12170 29469
rect 12130 29282 12182 29288
rect 55068 29282 55120 29288
rect 54967 29249 55068 29277
rect 12130 29224 12182 29230
rect 55068 29224 55120 29230
rect 12130 29042 12182 29048
rect 55068 29042 55120 29048
rect 54967 28995 55068 29023
rect 12130 28984 12182 28990
rect 55068 28984 55120 28990
rect 12142 28803 12170 28984
rect 12142 28775 12283 28803
rect 12142 28679 12283 28707
rect 12142 28498 12170 28679
rect 12130 28492 12182 28498
rect 55068 28492 55120 28498
rect 54967 28459 55068 28487
rect 12130 28434 12182 28440
rect 55068 28434 55120 28440
rect 12130 28252 12182 28258
rect 55068 28252 55120 28258
rect 54967 28205 55068 28233
rect 12130 28194 12182 28200
rect 55068 28194 55120 28200
rect 12142 28013 12170 28194
rect 12142 27985 12283 28013
rect 12142 27889 12283 27917
rect 12142 27708 12170 27889
rect 12130 27702 12182 27708
rect 55068 27702 55120 27708
rect 54967 27669 55068 27697
rect 12130 27644 12182 27650
rect 55068 27644 55120 27650
rect 12130 27462 12182 27468
rect 55068 27462 55120 27468
rect 54967 27415 55068 27443
rect 12130 27404 12182 27410
rect 55068 27404 55120 27410
rect 12142 27223 12170 27404
rect 12142 27195 12283 27223
rect 12142 27099 12283 27127
rect 12142 26918 12170 27099
rect 12130 26912 12182 26918
rect 55068 26912 55120 26918
rect 54967 26879 55068 26907
rect 12130 26854 12182 26860
rect 55068 26854 55120 26860
rect 12130 26672 12182 26678
rect 55068 26672 55120 26678
rect 54967 26625 55068 26653
rect 12130 26614 12182 26620
rect 55068 26614 55120 26620
rect 12142 26433 12170 26614
rect 12142 26405 12283 26433
rect 12142 26309 12283 26337
rect 12142 26128 12170 26309
rect 12130 26122 12182 26128
rect 55068 26122 55120 26128
rect 54967 26089 55068 26117
rect 12130 26064 12182 26070
rect 55068 26064 55120 26070
rect 12130 25882 12182 25888
rect 55068 25882 55120 25888
rect 54967 25835 55068 25863
rect 12130 25824 12182 25830
rect 55068 25824 55120 25830
rect 12142 25643 12170 25824
rect 12142 25615 12283 25643
rect 12142 25519 12283 25547
rect 12142 25338 12170 25519
rect 12130 25332 12182 25338
rect 55068 25332 55120 25338
rect 54967 25299 55068 25327
rect 12130 25274 12182 25280
rect 55068 25274 55120 25280
rect 12130 25092 12182 25098
rect 55068 25092 55120 25098
rect 54967 25045 55068 25073
rect 12130 25034 12182 25040
rect 55068 25034 55120 25040
rect 12142 24853 12170 25034
rect 12142 24825 12283 24853
rect 12142 24729 12283 24757
rect 12142 24548 12170 24729
rect 12130 24542 12182 24548
rect 55068 24542 55120 24548
rect 54967 24509 55068 24537
rect 12130 24484 12182 24490
rect 55068 24484 55120 24490
rect 12130 24302 12182 24308
rect 55068 24302 55120 24308
rect 54967 24255 55068 24283
rect 12130 24244 12182 24250
rect 55068 24244 55120 24250
rect 12142 24063 12170 24244
rect 12142 24035 12283 24063
rect 12142 23939 12283 23967
rect 12142 23758 12170 23939
rect 12130 23752 12182 23758
rect 55068 23752 55120 23758
rect 54967 23719 55068 23747
rect 12130 23694 12182 23700
rect 55068 23694 55120 23700
rect 12130 23512 12182 23518
rect 55068 23512 55120 23518
rect 54967 23465 55068 23493
rect 12130 23454 12182 23460
rect 55068 23454 55120 23460
rect 12142 23273 12170 23454
rect 12142 23245 12283 23273
rect 12142 23149 12283 23177
rect 12142 22968 12170 23149
rect 12130 22962 12182 22968
rect 55068 22962 55120 22968
rect 54967 22929 55068 22957
rect 12130 22904 12182 22910
rect 55068 22904 55120 22910
rect 12130 22722 12182 22728
rect 55068 22722 55120 22728
rect 54967 22675 55068 22703
rect 12130 22664 12182 22670
rect 55068 22664 55120 22670
rect 12142 22483 12170 22664
rect 12142 22455 12283 22483
rect 12142 22359 12283 22387
rect 12142 22178 12170 22359
rect 12130 22172 12182 22178
rect 55068 22172 55120 22178
rect 54967 22139 55068 22167
rect 12130 22114 12182 22120
rect 55068 22114 55120 22120
rect 12130 21932 12182 21938
rect 55068 21932 55120 21938
rect 54967 21885 55068 21913
rect 12130 21874 12182 21880
rect 55068 21874 55120 21880
rect 12142 21693 12170 21874
rect 12142 21665 12283 21693
rect 12142 21569 12283 21597
rect 12142 21388 12170 21569
rect 12130 21382 12182 21388
rect 55068 21382 55120 21388
rect 54967 21349 55068 21377
rect 12130 21324 12182 21330
rect 55068 21324 55120 21330
rect 12130 21142 12182 21148
rect 55068 21142 55120 21148
rect 54967 21095 55068 21123
rect 12130 21084 12182 21090
rect 55068 21084 55120 21090
rect 12142 20903 12170 21084
rect 12142 20875 12283 20903
rect 12142 20779 12283 20807
rect 12142 20598 12170 20779
rect 12130 20592 12182 20598
rect 55068 20592 55120 20598
rect 54967 20559 55068 20587
rect 12130 20534 12182 20540
rect 55068 20534 55120 20540
rect 12130 20352 12182 20358
rect 55068 20352 55120 20358
rect 54967 20305 55068 20333
rect 12130 20294 12182 20300
rect 55068 20294 55120 20300
rect 12142 20113 12170 20294
rect 12142 20085 12283 20113
rect 12142 19989 12283 20017
rect 12142 19808 12170 19989
rect 12130 19802 12182 19808
rect 55068 19802 55120 19808
rect 54967 19769 55068 19797
rect 12130 19744 12182 19750
rect 55068 19744 55120 19750
rect 12130 19562 12182 19568
rect 55068 19562 55120 19568
rect 54967 19515 55068 19543
rect 12130 19504 12182 19510
rect 55068 19504 55120 19510
rect 12142 19323 12170 19504
rect 12142 19295 12283 19323
rect 12142 19199 12283 19227
rect 12142 19018 12170 19199
rect 12130 19012 12182 19018
rect 55068 19012 55120 19018
rect 54967 18979 55068 19007
rect 12130 18954 12182 18960
rect 55068 18954 55120 18960
rect 12130 18772 12182 18778
rect 55068 18772 55120 18778
rect 54967 18725 55068 18753
rect 12130 18714 12182 18720
rect 55068 18714 55120 18720
rect 12142 18533 12170 18714
rect 12142 18505 12283 18533
rect 12142 18409 12283 18437
rect 12142 18228 12170 18409
rect 12130 18222 12182 18228
rect 55068 18222 55120 18228
rect 54967 18189 55068 18217
rect 12130 18164 12182 18170
rect 55068 18164 55120 18170
rect 12130 17982 12182 17988
rect 55068 17982 55120 17988
rect 54967 17935 55068 17963
rect 12130 17924 12182 17930
rect 55068 17924 55120 17930
rect 12142 17743 12170 17924
rect 12142 17715 12283 17743
rect 12142 17619 12283 17647
rect 12142 17438 12170 17619
rect 12130 17432 12182 17438
rect 55068 17432 55120 17438
rect 54967 17399 55068 17427
rect 12130 17374 12182 17380
rect 55068 17374 55120 17380
rect 12130 17192 12182 17198
rect 55068 17192 55120 17198
rect 54967 17145 55068 17173
rect 12130 17134 12182 17140
rect 55068 17134 55120 17140
rect 12142 16953 12170 17134
rect 12142 16925 12283 16953
rect 12142 16829 12283 16857
rect 12142 16648 12170 16829
rect 12130 16642 12182 16648
rect 55068 16642 55120 16648
rect 54967 16609 55068 16637
rect 12130 16584 12182 16590
rect 55068 16584 55120 16590
rect 12130 16402 12182 16408
rect 55068 16402 55120 16408
rect 54967 16355 55068 16383
rect 12130 16344 12182 16350
rect 55068 16344 55120 16350
rect 12142 16163 12170 16344
rect 12142 16135 12283 16163
rect 12142 16039 12283 16067
rect 12142 15858 12170 16039
rect 12130 15852 12182 15858
rect 55068 15852 55120 15858
rect 54967 15819 55068 15847
rect 12130 15794 12182 15800
rect 55068 15794 55120 15800
rect 12130 15612 12182 15618
rect 55068 15612 55120 15618
rect 54967 15565 55068 15593
rect 12130 15554 12182 15560
rect 55068 15554 55120 15560
rect 12142 15373 12170 15554
rect 12142 15345 12283 15373
rect 12142 15249 12283 15277
rect 12142 15068 12170 15249
rect 12130 15062 12182 15068
rect 55068 15062 55120 15068
rect 54967 15029 55068 15057
rect 12130 15004 12182 15010
rect 55068 15004 55120 15010
rect 12130 14822 12182 14828
rect 55068 14822 55120 14828
rect 54967 14775 55068 14803
rect 12130 14764 12182 14770
rect 55068 14764 55120 14770
rect 12142 14583 12170 14764
rect 12142 14555 12283 14583
rect 12142 14459 12283 14487
rect 12142 14278 12170 14459
rect 12130 14272 12182 14278
rect 55068 14272 55120 14278
rect 54967 14239 55068 14267
rect 12130 14214 12182 14220
rect 55068 14214 55120 14220
rect 12130 14032 12182 14038
rect 55068 14032 55120 14038
rect 54967 13985 55068 14013
rect 12130 13974 12182 13980
rect 55068 13974 55120 13980
rect 12142 13793 12170 13974
rect 12142 13765 12283 13793
rect 12142 13669 12283 13697
rect 12142 13488 12170 13669
rect 12130 13482 12182 13488
rect 55068 13482 55120 13488
rect 54967 13449 55068 13477
rect 12130 13424 12182 13430
rect 55068 13424 55120 13430
rect 12130 13242 12182 13248
rect 55068 13242 55120 13248
rect 54967 13195 55068 13223
rect 12130 13184 12182 13190
rect 55068 13184 55120 13190
rect 12142 13003 12170 13184
rect 12142 12975 12283 13003
rect 12142 12879 12283 12907
rect 12142 12698 12170 12879
rect 12130 12692 12182 12698
rect 55068 12692 55120 12698
rect 54967 12659 55068 12687
rect 12130 12634 12182 12640
rect 55068 12634 55120 12640
rect 12130 12452 12182 12458
rect 55068 12452 55120 12458
rect 54967 12405 55068 12433
rect 12130 12394 12182 12400
rect 55068 12394 55120 12400
rect 12142 12213 12170 12394
rect 12142 12185 12283 12213
rect 12142 12089 12283 12117
rect 12142 11908 12170 12089
rect 12130 11902 12182 11908
rect 55068 11902 55120 11908
rect 54967 11869 55068 11897
rect 12130 11844 12182 11850
rect 55068 11844 55120 11850
rect 12130 11662 12182 11668
rect 55068 11662 55120 11668
rect 54967 11615 55068 11643
rect 12130 11604 12182 11610
rect 55068 11604 55120 11610
rect 12142 11423 12170 11604
rect 12142 11395 12283 11423
rect 12142 11299 12283 11327
rect 12142 11118 12170 11299
rect 12130 11112 12182 11118
rect 55068 11112 55120 11118
rect 54967 11079 55068 11107
rect 12130 11054 12182 11060
rect 55068 11054 55120 11060
rect 12130 10872 12182 10878
rect 55068 10872 55120 10878
rect 54967 10825 55068 10853
rect 12130 10814 12182 10820
rect 55068 10814 55120 10820
rect 12142 10633 12170 10814
rect 12142 10605 12283 10633
rect 12142 10509 12283 10537
rect 12142 10328 12170 10509
rect 12130 10322 12182 10328
rect 55068 10322 55120 10328
rect 54967 10289 55068 10317
rect 12130 10264 12182 10270
rect 55068 10264 55120 10270
rect 12130 10082 12182 10088
rect 12130 10024 12182 10030
rect 7960 9863 7988 9891
rect 12142 9843 12170 10024
rect 12142 9815 12283 9843
rect 11663 8442 11691 9386
rect 11649 8433 11705 8442
rect 11649 8368 11705 8377
rect 6729 7663 6785 7672
rect 6729 7598 6785 7607
rect 7128 6956 7184 6965
rect 7128 6891 7184 6900
rect 7757 6956 7813 6965
rect 7757 6891 7813 6900
rect 7771 6755 7799 6891
rect 7757 6746 7813 6755
rect 7757 6681 7813 6690
rect 7621 6622 7677 6631
rect 7621 6557 7677 6566
rect 6729 6249 6785 6258
rect 6729 6184 6785 6193
rect 7635 5551 7663 6557
rect 7128 5542 7184 5551
rect 7128 5477 7184 5486
rect 7621 5542 7677 5551
rect 7621 5477 7677 5486
rect 6729 4835 6785 4844
rect 6729 4770 6785 4779
rect 11663 49 11691 8368
rect 11787 5915 11815 9386
rect 11773 5906 11829 5915
rect 11773 5841 11829 5850
rect 11787 49 11815 5841
rect 11911 604 11939 9386
rect 13549 8284 13605 8293
rect 13549 8219 13605 8228
rect 11897 595 11953 604
rect 11897 530 11953 539
rect 11911 49 11939 530
rect 13643 305 13671 333
rect 23627 305 23655 333
rect 33611 305 33639 333
rect 43595 305 43623 333
<< via2 >>
rect 55263 65006 55319 65062
rect 53645 62682 53701 62684
rect 53645 62630 53647 62682
rect 53647 62630 53699 62682
rect 53699 62630 53701 62682
rect 53645 62628 53701 62630
rect 60341 66131 60397 66133
rect 60341 66079 60343 66131
rect 60343 66079 60395 66131
rect 60395 66079 60397 66131
rect 60341 66077 60397 66079
rect 59337 65370 59393 65426
rect 59942 65424 59998 65426
rect 59942 65372 59944 65424
rect 59944 65372 59996 65424
rect 59996 65372 59998 65424
rect 59942 65370 59998 65372
rect 60341 64717 60397 64719
rect 60341 64665 60343 64717
rect 60343 64665 60395 64717
rect 60395 64665 60397 64717
rect 60341 64663 60397 64665
rect 59337 64290 59393 64346
rect 59201 64166 59257 64222
rect 59201 63956 59257 64012
rect 59942 64010 59998 64012
rect 59942 63958 59944 64010
rect 59944 63958 59996 64010
rect 59996 63958 59998 64010
rect 59942 63956 59998 63958
rect 60341 63303 60397 63305
rect 60341 63251 60343 63303
rect 60343 63251 60395 63303
rect 60395 63251 60397 63303
rect 60341 63249 60397 63251
rect 55387 62479 55443 62535
rect 11649 8377 11705 8433
rect 6729 7661 6785 7663
rect 6729 7609 6731 7661
rect 6731 7609 6783 7661
rect 6783 7609 6785 7661
rect 6729 7607 6785 7609
rect 7128 6954 7184 6956
rect 7128 6902 7130 6954
rect 7130 6902 7182 6954
rect 7182 6902 7184 6954
rect 7128 6900 7184 6902
rect 7757 6900 7813 6956
rect 7757 6690 7813 6746
rect 7621 6566 7677 6622
rect 6729 6247 6785 6249
rect 6729 6195 6731 6247
rect 6731 6195 6783 6247
rect 6783 6195 6785 6247
rect 6729 6193 6785 6195
rect 7128 5540 7184 5542
rect 7128 5488 7130 5540
rect 7130 5488 7182 5540
rect 7182 5488 7184 5540
rect 7128 5486 7184 5488
rect 7621 5486 7677 5542
rect 6729 4833 6785 4835
rect 6729 4781 6731 4833
rect 6731 4781 6783 4833
rect 6783 4781 6785 4833
rect 6729 4779 6785 4781
rect 11773 5850 11829 5906
rect 13549 8282 13605 8284
rect 13549 8230 13551 8282
rect 13551 8230 13603 8282
rect 13603 8230 13605 8282
rect 13549 8228 13605 8230
rect 11897 539 11953 595
<< metal3 >>
rect 13989 67071 14087 67169
rect 15237 67071 15335 67169
rect 16485 67071 16583 67169
rect 17733 67071 17831 67169
rect 18981 67071 19079 67169
rect 20229 67071 20327 67169
rect 21477 67071 21575 67169
rect 22725 67071 22823 67169
rect 23973 67071 24071 67169
rect 25221 67071 25319 67169
rect 26469 67071 26567 67169
rect 27717 67071 27815 67169
rect 28965 67071 29063 67169
rect 30213 67071 30311 67169
rect 31461 67071 31559 67169
rect 32709 67071 32807 67169
rect 33957 67071 34055 67169
rect 35205 67071 35303 67169
rect 36453 67071 36551 67169
rect 37701 67071 37799 67169
rect 38949 67071 39047 67169
rect 40197 67071 40295 67169
rect 41445 67071 41543 67169
rect 42693 67071 42791 67169
rect 43941 67071 44039 67169
rect 45189 67071 45287 67169
rect 46437 67071 46535 67169
rect 47685 67071 47783 67169
rect 48933 67071 49031 67169
rect 50181 67071 50279 67169
rect 51429 67071 51527 67169
rect 52677 67071 52775 67169
rect 13989 66749 14087 66847
rect 15237 66749 15335 66847
rect 16485 66749 16583 66847
rect 17733 66749 17831 66847
rect 18981 66749 19079 66847
rect 20229 66749 20327 66847
rect 21477 66749 21575 66847
rect 22725 66749 22823 66847
rect 23973 66749 24071 66847
rect 25221 66749 25319 66847
rect 26469 66749 26567 66847
rect 27717 66749 27815 66847
rect 28965 66749 29063 66847
rect 30213 66749 30311 66847
rect 31461 66749 31559 66847
rect 32709 66749 32807 66847
rect 33957 66749 34055 66847
rect 35205 66749 35303 66847
rect 36453 66749 36551 66847
rect 37701 66749 37799 66847
rect 38949 66749 39047 66847
rect 40197 66749 40295 66847
rect 41445 66749 41543 66847
rect 42693 66749 42791 66847
rect 43941 66749 44039 66847
rect 45189 66749 45287 66847
rect 46437 66749 46535 66847
rect 47685 66749 47783 66847
rect 48933 66749 49031 66847
rect 50181 66749 50279 66847
rect 51429 66749 51527 66847
rect 52677 66749 52775 66847
rect 60320 66133 60418 66154
rect 60320 66077 60341 66133
rect 60397 66077 60418 66133
rect 60320 66056 60418 66077
rect 13977 65911 14075 66009
rect 15225 65911 15323 66009
rect 16473 65911 16571 66009
rect 17721 65911 17819 66009
rect 18969 65911 19067 66009
rect 20217 65911 20315 66009
rect 21465 65911 21563 66009
rect 22713 65911 22811 66009
rect 23961 65911 24059 66009
rect 25209 65911 25307 66009
rect 26457 65911 26555 66009
rect 27705 65911 27803 66009
rect 28953 65911 29051 66009
rect 30201 65911 30299 66009
rect 31449 65911 31547 66009
rect 32697 65911 32795 66009
rect 33945 65911 34043 66009
rect 35193 65911 35291 66009
rect 36441 65911 36539 66009
rect 37689 65911 37787 66009
rect 38937 65911 39035 66009
rect 40185 65911 40283 66009
rect 41433 65911 41531 66009
rect 42681 65911 42779 66009
rect 43929 65911 44027 66009
rect 45177 65911 45275 66009
rect 46425 65911 46523 66009
rect 47673 65911 47771 66009
rect 48921 65911 49019 66009
rect 50169 65911 50267 66009
rect 51417 65911 51515 66009
rect 52665 65911 52763 66009
rect 59332 65428 59398 65431
rect 59937 65428 60003 65431
rect 59332 65426 60003 65428
rect 59332 65370 59337 65426
rect 59393 65370 59942 65426
rect 59998 65370 60003 65426
rect 59332 65368 60003 65370
rect 59332 65365 59398 65368
rect 59937 65365 60003 65368
rect 14059 65137 14157 65235
rect 15307 65137 15405 65235
rect 16555 65137 16653 65235
rect 17803 65137 17901 65235
rect 19051 65137 19149 65235
rect 20299 65137 20397 65235
rect 21547 65137 21645 65235
rect 22795 65137 22893 65235
rect 24043 65137 24141 65235
rect 25291 65137 25389 65235
rect 26539 65137 26637 65235
rect 27787 65137 27885 65235
rect 29035 65137 29133 65235
rect 30283 65137 30381 65235
rect 31531 65137 31629 65235
rect 32779 65137 32877 65235
rect 34027 65137 34125 65235
rect 35275 65137 35373 65235
rect 36523 65137 36621 65235
rect 37771 65137 37869 65235
rect 39019 65137 39117 65235
rect 40267 65137 40365 65235
rect 41515 65137 41613 65235
rect 42763 65137 42861 65235
rect 44011 65137 44109 65235
rect 45259 65137 45357 65235
rect 46507 65137 46605 65235
rect 47755 65137 47853 65235
rect 49003 65137 49101 65235
rect 50251 65137 50349 65235
rect 51499 65137 51597 65235
rect 52747 65137 52845 65235
rect 55258 65064 55324 65067
rect 32564 65062 55324 65064
rect 32564 65006 55263 65062
rect 55319 65006 55324 65062
rect 32564 65004 55324 65006
rect 55258 65001 55324 65004
rect 60320 64719 60418 64740
rect 60320 64663 60341 64719
rect 60397 64663 60418 64719
rect 60320 64642 60418 64663
rect 59332 64348 59398 64351
rect 53563 64346 59398 64348
rect 53563 64290 59337 64346
rect 59393 64290 59398 64346
rect 53563 64288 59398 64290
rect 59332 64285 59398 64288
rect 59196 64224 59262 64227
rect 53563 64222 59262 64224
rect 53563 64166 59201 64222
rect 59257 64166 59262 64222
rect 53563 64164 59262 64166
rect 59196 64161 59262 64164
rect 59196 64014 59262 64017
rect 59937 64014 60003 64017
rect 59196 64012 60003 64014
rect 59196 63956 59201 64012
rect 59257 63956 59942 64012
rect 59998 63956 60003 64012
rect 59196 63954 60003 63956
rect 59196 63951 59262 63954
rect 59937 63951 60003 63954
rect 14232 63388 14330 63486
rect 15480 63388 15578 63486
rect 16728 63388 16826 63486
rect 17976 63388 18074 63486
rect 19224 63388 19322 63486
rect 20472 63388 20570 63486
rect 21720 63388 21818 63486
rect 22968 63388 23066 63486
rect 24216 63388 24314 63486
rect 25464 63388 25562 63486
rect 26712 63388 26810 63486
rect 27960 63388 28058 63486
rect 29208 63388 29306 63486
rect 30456 63388 30554 63486
rect 31704 63388 31802 63486
rect 32952 63388 33050 63486
rect 34200 63388 34298 63486
rect 35448 63388 35546 63486
rect 36696 63388 36794 63486
rect 37944 63388 38042 63486
rect 39192 63388 39290 63486
rect 40440 63388 40538 63486
rect 41688 63388 41786 63486
rect 42936 63388 43034 63486
rect 44184 63388 44282 63486
rect 45432 63388 45530 63486
rect 46680 63388 46778 63486
rect 47928 63388 48026 63486
rect 49176 63388 49274 63486
rect 50424 63388 50522 63486
rect 51672 63388 51770 63486
rect 52920 63388 53018 63486
rect 60320 63305 60418 63326
rect 60320 63249 60341 63305
rect 60397 63249 60418 63305
rect 60320 63228 60418 63249
rect 53640 62686 53706 62689
rect 53640 62684 67334 62686
rect 53640 62628 53645 62684
rect 53701 62628 67334 62684
rect 53640 62626 67334 62628
rect 53640 62623 53706 62626
rect 55382 62537 55448 62540
rect 33250 62535 55448 62537
rect 33250 62479 55387 62535
rect 55443 62479 55448 62535
rect 33250 62477 55448 62479
rect 55382 62474 55448 62477
rect 13801 61839 13899 61937
rect 14663 61839 14761 61937
rect 15049 61839 15147 61937
rect 15911 61839 16009 61937
rect 16297 61839 16395 61937
rect 17159 61839 17257 61937
rect 17545 61839 17643 61937
rect 18407 61839 18505 61937
rect 18793 61839 18891 61937
rect 19655 61839 19753 61937
rect 20041 61839 20139 61937
rect 20903 61839 21001 61937
rect 21289 61839 21387 61937
rect 22151 61839 22249 61937
rect 22537 61839 22635 61937
rect 23399 61839 23497 61937
rect 23785 61839 23883 61937
rect 24647 61839 24745 61937
rect 25033 61839 25131 61937
rect 25895 61839 25993 61937
rect 26281 61839 26379 61937
rect 27143 61839 27241 61937
rect 27529 61839 27627 61937
rect 28391 61839 28489 61937
rect 28777 61839 28875 61937
rect 29639 61839 29737 61937
rect 30025 61839 30123 61937
rect 30887 61839 30985 61937
rect 31273 61839 31371 61937
rect 32135 61839 32233 61937
rect 32521 61839 32619 61937
rect 33383 61839 33481 61937
rect 33769 61839 33867 61937
rect 34631 61839 34729 61937
rect 35017 61839 35115 61937
rect 35879 61839 35977 61937
rect 36265 61839 36363 61937
rect 37127 61839 37225 61937
rect 37513 61839 37611 61937
rect 38375 61839 38473 61937
rect 38761 61839 38859 61937
rect 39623 61839 39721 61937
rect 40009 61839 40107 61937
rect 40871 61839 40969 61937
rect 41257 61839 41355 61937
rect 42119 61839 42217 61937
rect 42505 61839 42603 61937
rect 43367 61839 43465 61937
rect 43753 61839 43851 61937
rect 44615 61839 44713 61937
rect 45001 61839 45099 61937
rect 45863 61839 45961 61937
rect 46249 61839 46347 61937
rect 47111 61839 47209 61937
rect 47497 61839 47595 61937
rect 48359 61839 48457 61937
rect 48745 61839 48843 61937
rect 49607 61839 49705 61937
rect 49993 61839 50091 61937
rect 50855 61839 50953 61937
rect 51241 61839 51339 61937
rect 52103 61839 52201 61937
rect 52489 61839 52587 61937
rect 53351 61839 53449 61937
rect 53737 61839 53835 61937
rect 13296 61248 13394 61346
rect 13920 61248 14018 61346
rect 14544 61248 14642 61346
rect 15168 61248 15266 61346
rect 15792 61248 15890 61346
rect 16416 61248 16514 61346
rect 17040 61248 17138 61346
rect 17664 61248 17762 61346
rect 18288 61248 18386 61346
rect 18912 61248 19010 61346
rect 19536 61248 19634 61346
rect 20160 61248 20258 61346
rect 20784 61248 20882 61346
rect 21408 61248 21506 61346
rect 22032 61248 22130 61346
rect 22656 61248 22754 61346
rect 23280 61248 23378 61346
rect 23904 61248 24002 61346
rect 24528 61248 24626 61346
rect 25152 61248 25250 61346
rect 25776 61248 25874 61346
rect 26400 61248 26498 61346
rect 27024 61248 27122 61346
rect 27648 61248 27746 61346
rect 28272 61248 28370 61346
rect 28896 61248 28994 61346
rect 29520 61248 29618 61346
rect 30144 61248 30242 61346
rect 30768 61248 30866 61346
rect 31392 61248 31490 61346
rect 32016 61248 32114 61346
rect 32640 61248 32738 61346
rect 33264 61248 33362 61346
rect 33888 61248 33986 61346
rect 34512 61248 34610 61346
rect 35136 61248 35234 61346
rect 35760 61248 35858 61346
rect 36384 61248 36482 61346
rect 37008 61248 37106 61346
rect 37632 61248 37730 61346
rect 38256 61248 38354 61346
rect 38880 61248 38978 61346
rect 39504 61248 39602 61346
rect 40128 61248 40226 61346
rect 40752 61248 40850 61346
rect 41376 61248 41474 61346
rect 42000 61248 42098 61346
rect 42624 61248 42722 61346
rect 43248 61248 43346 61346
rect 43872 61248 43970 61346
rect 44496 61248 44594 61346
rect 45120 61248 45218 61346
rect 45744 61248 45842 61346
rect 46368 61248 46466 61346
rect 46992 61248 47090 61346
rect 47616 61248 47714 61346
rect 48240 61248 48338 61346
rect 48864 61248 48962 61346
rect 49488 61248 49586 61346
rect 50112 61248 50210 61346
rect 50736 61248 50834 61346
rect 51360 61248 51458 61346
rect 51984 61248 52082 61346
rect 52608 61248 52706 61346
rect 53232 61248 53330 61346
rect 53856 61248 53954 61346
rect 12234 61034 12332 61132
rect 54918 61034 55016 61132
rect 55944 60884 56042 60982
rect 58635 60872 58733 60970
rect 59467 60878 59565 60976
rect 12600 60687 12698 60785
rect 54552 60687 54650 60785
rect 12600 60450 12698 60548
rect 54552 60450 54650 60548
rect 6025 60315 6123 60413
rect 6450 60315 6548 60413
rect 6882 60315 6980 60413
rect 7264 60292 7362 60390
rect 7660 60292 7758 60390
rect 59492 60292 59590 60390
rect 59888 60292 59986 60390
rect 60270 60315 60368 60413
rect 60702 60315 60800 60413
rect 61127 60315 61225 60413
rect 12600 60134 12698 60232
rect 54552 60134 54650 60232
rect 6025 59941 6123 60039
rect 6450 59883 6548 59981
rect 6882 59883 6980 59981
rect 7264 59897 7362 59995
rect 7660 59897 7758 59995
rect 12600 59897 12698 59995
rect 54552 59897 54650 59995
rect 59492 59897 59590 59995
rect 59888 59897 59986 59995
rect 60270 59883 60368 59981
rect 60702 59883 60800 59981
rect 61127 59941 61225 60039
rect 12600 59660 12698 59758
rect 54552 59660 54650 59758
rect 6025 59525 6123 59623
rect 6450 59525 6548 59623
rect 6882 59525 6980 59623
rect 7264 59502 7362 59600
rect 7660 59502 7758 59600
rect 59492 59502 59590 59600
rect 59888 59502 59986 59600
rect 60270 59525 60368 59623
rect 60702 59525 60800 59623
rect 61127 59525 61225 59623
rect 12600 59344 12698 59442
rect 54552 59344 54650 59442
rect 6025 59151 6123 59249
rect 6450 59093 6548 59191
rect 6882 59093 6980 59191
rect 7264 59107 7362 59205
rect 7660 59107 7758 59205
rect 12600 59107 12698 59205
rect 54552 59107 54650 59205
rect 59492 59107 59590 59205
rect 59888 59107 59986 59205
rect 60270 59093 60368 59191
rect 60702 59093 60800 59191
rect 61127 59151 61225 59249
rect 12600 58870 12698 58968
rect 54552 58870 54650 58968
rect 6025 58735 6123 58833
rect 6450 58735 6548 58833
rect 6882 58735 6980 58833
rect 7264 58712 7362 58810
rect 7660 58712 7758 58810
rect 59492 58712 59590 58810
rect 59888 58712 59986 58810
rect 60270 58735 60368 58833
rect 60702 58735 60800 58833
rect 61127 58735 61225 58833
rect 12600 58554 12698 58652
rect 54552 58554 54650 58652
rect 6025 58361 6123 58459
rect 6450 58303 6548 58401
rect 6882 58303 6980 58401
rect 7264 58317 7362 58415
rect 7660 58317 7758 58415
rect 12600 58317 12698 58415
rect 54552 58317 54650 58415
rect 59492 58317 59590 58415
rect 59888 58317 59986 58415
rect 60270 58303 60368 58401
rect 60702 58303 60800 58401
rect 61127 58361 61225 58459
rect 12600 58080 12698 58178
rect 54552 58080 54650 58178
rect 6025 57945 6123 58043
rect 6450 57945 6548 58043
rect 6882 57945 6980 58043
rect 7264 57922 7362 58020
rect 7660 57922 7758 58020
rect 59492 57922 59590 58020
rect 59888 57922 59986 58020
rect 60270 57945 60368 58043
rect 60702 57945 60800 58043
rect 61127 57945 61225 58043
rect 12600 57764 12698 57862
rect 54552 57764 54650 57862
rect 6025 57571 6123 57669
rect 6450 57513 6548 57611
rect 6882 57513 6980 57611
rect 7264 57527 7362 57625
rect 7660 57527 7758 57625
rect 12600 57527 12698 57625
rect 54552 57527 54650 57625
rect 59492 57527 59590 57625
rect 59888 57527 59986 57625
rect 60270 57513 60368 57611
rect 60702 57513 60800 57611
rect 61127 57571 61225 57669
rect 12600 57290 12698 57388
rect 54552 57290 54650 57388
rect 6025 57155 6123 57253
rect 6450 57155 6548 57253
rect 6882 57155 6980 57253
rect 7264 57132 7362 57230
rect 7660 57132 7758 57230
rect 59492 57132 59590 57230
rect 59888 57132 59986 57230
rect 60270 57155 60368 57253
rect 60702 57155 60800 57253
rect 61127 57155 61225 57253
rect 12600 56974 12698 57072
rect 54552 56974 54650 57072
rect 6025 56781 6123 56879
rect 6450 56723 6548 56821
rect 6882 56723 6980 56821
rect 7264 56737 7362 56835
rect 7660 56737 7758 56835
rect 12600 56737 12698 56835
rect 54552 56737 54650 56835
rect 59492 56737 59590 56835
rect 59888 56737 59986 56835
rect 60270 56723 60368 56821
rect 60702 56723 60800 56821
rect 61127 56781 61225 56879
rect 12600 56500 12698 56598
rect 54552 56500 54650 56598
rect 6025 56365 6123 56463
rect 6450 56365 6548 56463
rect 6882 56365 6980 56463
rect 7264 56342 7362 56440
rect 7660 56342 7758 56440
rect 59492 56342 59590 56440
rect 59888 56342 59986 56440
rect 60270 56365 60368 56463
rect 60702 56365 60800 56463
rect 61127 56365 61225 56463
rect 12600 56184 12698 56282
rect 54552 56184 54650 56282
rect 6025 55991 6123 56089
rect 6450 55933 6548 56031
rect 6882 55933 6980 56031
rect 7264 55947 7362 56045
rect 7660 55947 7758 56045
rect 12600 55947 12698 56045
rect 54552 55947 54650 56045
rect 59492 55947 59590 56045
rect 59888 55947 59986 56045
rect 60270 55933 60368 56031
rect 60702 55933 60800 56031
rect 61127 55991 61225 56089
rect 12600 55710 12698 55808
rect 54552 55710 54650 55808
rect 6025 55575 6123 55673
rect 6450 55575 6548 55673
rect 6882 55575 6980 55673
rect 7264 55552 7362 55650
rect 7660 55552 7758 55650
rect 59492 55552 59590 55650
rect 59888 55552 59986 55650
rect 60270 55575 60368 55673
rect 60702 55575 60800 55673
rect 61127 55575 61225 55673
rect 12600 55394 12698 55492
rect 54552 55394 54650 55492
rect 6025 55201 6123 55299
rect 6450 55143 6548 55241
rect 6882 55143 6980 55241
rect 7264 55157 7362 55255
rect 7660 55157 7758 55255
rect 12600 55157 12698 55255
rect 54552 55157 54650 55255
rect 59492 55157 59590 55255
rect 59888 55157 59986 55255
rect 60270 55143 60368 55241
rect 60702 55143 60800 55241
rect 61127 55201 61225 55299
rect 12600 54920 12698 55018
rect 54552 54920 54650 55018
rect 6025 54785 6123 54883
rect 6450 54785 6548 54883
rect 6882 54785 6980 54883
rect 7264 54762 7362 54860
rect 7660 54762 7758 54860
rect 59492 54762 59590 54860
rect 59888 54762 59986 54860
rect 60270 54785 60368 54883
rect 60702 54785 60800 54883
rect 61127 54785 61225 54883
rect 12600 54604 12698 54702
rect 54552 54604 54650 54702
rect 6025 54411 6123 54509
rect 6450 54353 6548 54451
rect 6882 54353 6980 54451
rect 7264 54367 7362 54465
rect 7660 54367 7758 54465
rect 12600 54367 12698 54465
rect 54552 54367 54650 54465
rect 59492 54367 59590 54465
rect 59888 54367 59986 54465
rect 60270 54353 60368 54451
rect 60702 54353 60800 54451
rect 61127 54411 61225 54509
rect 12600 54130 12698 54228
rect 54552 54130 54650 54228
rect 6025 53995 6123 54093
rect 6450 53995 6548 54093
rect 6882 53995 6980 54093
rect 7264 53972 7362 54070
rect 7660 53972 7758 54070
rect 59492 53972 59590 54070
rect 59888 53972 59986 54070
rect 60270 53995 60368 54093
rect 60702 53995 60800 54093
rect 61127 53995 61225 54093
rect 12600 53814 12698 53912
rect 54552 53814 54650 53912
rect 6025 53621 6123 53719
rect 6450 53563 6548 53661
rect 6882 53563 6980 53661
rect 7264 53577 7362 53675
rect 7660 53577 7758 53675
rect 12600 53577 12698 53675
rect 54552 53577 54650 53675
rect 59492 53577 59590 53675
rect 59888 53577 59986 53675
rect 60270 53563 60368 53661
rect 60702 53563 60800 53661
rect 61127 53621 61225 53719
rect 12600 53340 12698 53438
rect 54552 53340 54650 53438
rect 6025 53205 6123 53303
rect 6450 53205 6548 53303
rect 6882 53205 6980 53303
rect 7264 53182 7362 53280
rect 7660 53182 7758 53280
rect 59492 53182 59590 53280
rect 59888 53182 59986 53280
rect 60270 53205 60368 53303
rect 60702 53205 60800 53303
rect 61127 53205 61225 53303
rect 12600 53024 12698 53122
rect 54552 53024 54650 53122
rect 6025 52831 6123 52929
rect 6450 52773 6548 52871
rect 6882 52773 6980 52871
rect 7264 52787 7362 52885
rect 7660 52787 7758 52885
rect 12600 52787 12698 52885
rect 54552 52787 54650 52885
rect 59492 52787 59590 52885
rect 59888 52787 59986 52885
rect 60270 52773 60368 52871
rect 60702 52773 60800 52871
rect 61127 52831 61225 52929
rect 12600 52550 12698 52648
rect 54552 52550 54650 52648
rect 6025 52415 6123 52513
rect 6450 52415 6548 52513
rect 6882 52415 6980 52513
rect 7264 52392 7362 52490
rect 7660 52392 7758 52490
rect 59492 52392 59590 52490
rect 59888 52392 59986 52490
rect 60270 52415 60368 52513
rect 60702 52415 60800 52513
rect 61127 52415 61225 52513
rect 12600 52234 12698 52332
rect 54552 52234 54650 52332
rect 6025 52041 6123 52139
rect 6450 51983 6548 52081
rect 6882 51983 6980 52081
rect 7264 51997 7362 52095
rect 7660 51997 7758 52095
rect 12600 51997 12698 52095
rect 54552 51997 54650 52095
rect 59492 51997 59590 52095
rect 59888 51997 59986 52095
rect 60270 51983 60368 52081
rect 60702 51983 60800 52081
rect 61127 52041 61225 52139
rect 12600 51760 12698 51858
rect 54552 51760 54650 51858
rect 6025 51625 6123 51723
rect 6450 51625 6548 51723
rect 6882 51625 6980 51723
rect 7264 51602 7362 51700
rect 7660 51602 7758 51700
rect 59492 51602 59590 51700
rect 59888 51602 59986 51700
rect 60270 51625 60368 51723
rect 60702 51625 60800 51723
rect 61127 51625 61225 51723
rect 12600 51444 12698 51542
rect 54552 51444 54650 51542
rect 6025 51251 6123 51349
rect 6450 51193 6548 51291
rect 6882 51193 6980 51291
rect 7264 51207 7362 51305
rect 7660 51207 7758 51305
rect 12600 51207 12698 51305
rect 54552 51207 54650 51305
rect 59492 51207 59590 51305
rect 59888 51207 59986 51305
rect 60270 51193 60368 51291
rect 60702 51193 60800 51291
rect 61127 51251 61225 51349
rect 12600 50970 12698 51068
rect 54552 50970 54650 51068
rect 6025 50835 6123 50933
rect 6450 50835 6548 50933
rect 6882 50835 6980 50933
rect 7264 50812 7362 50910
rect 7660 50812 7758 50910
rect 59492 50812 59590 50910
rect 59888 50812 59986 50910
rect 60270 50835 60368 50933
rect 60702 50835 60800 50933
rect 61127 50835 61225 50933
rect 12600 50654 12698 50752
rect 54552 50654 54650 50752
rect 6025 50461 6123 50559
rect 6450 50403 6548 50501
rect 6882 50403 6980 50501
rect 7264 50417 7362 50515
rect 7660 50417 7758 50515
rect 12600 50417 12698 50515
rect 54552 50417 54650 50515
rect 59492 50417 59590 50515
rect 59888 50417 59986 50515
rect 60270 50403 60368 50501
rect 60702 50403 60800 50501
rect 61127 50461 61225 50559
rect 12600 50180 12698 50278
rect 54552 50180 54650 50278
rect 6025 50045 6123 50143
rect 6450 50045 6548 50143
rect 6882 50045 6980 50143
rect 7264 50022 7362 50120
rect 7660 50022 7758 50120
rect 59492 50022 59590 50120
rect 59888 50022 59986 50120
rect 60270 50045 60368 50143
rect 60702 50045 60800 50143
rect 61127 50045 61225 50143
rect 12600 49864 12698 49962
rect 54552 49864 54650 49962
rect 6025 49671 6123 49769
rect 6450 49613 6548 49711
rect 6882 49613 6980 49711
rect 7264 49627 7362 49725
rect 7660 49627 7758 49725
rect 12600 49627 12698 49725
rect 54552 49627 54650 49725
rect 59492 49627 59590 49725
rect 59888 49627 59986 49725
rect 60270 49613 60368 49711
rect 60702 49613 60800 49711
rect 61127 49671 61225 49769
rect 12600 49390 12698 49488
rect 54552 49390 54650 49488
rect 6025 49255 6123 49353
rect 6450 49255 6548 49353
rect 6882 49255 6980 49353
rect 7264 49232 7362 49330
rect 7660 49232 7758 49330
rect 59492 49232 59590 49330
rect 59888 49232 59986 49330
rect 60270 49255 60368 49353
rect 60702 49255 60800 49353
rect 61127 49255 61225 49353
rect 12600 49074 12698 49172
rect 54552 49074 54650 49172
rect 6025 48881 6123 48979
rect 6450 48823 6548 48921
rect 6882 48823 6980 48921
rect 7264 48837 7362 48935
rect 7660 48837 7758 48935
rect 12600 48837 12698 48935
rect 54552 48837 54650 48935
rect 59492 48837 59590 48935
rect 59888 48837 59986 48935
rect 60270 48823 60368 48921
rect 60702 48823 60800 48921
rect 61127 48881 61225 48979
rect 12600 48600 12698 48698
rect 54552 48600 54650 48698
rect 6025 48465 6123 48563
rect 6450 48465 6548 48563
rect 6882 48465 6980 48563
rect 7264 48442 7362 48540
rect 7660 48442 7758 48540
rect 59492 48442 59590 48540
rect 59888 48442 59986 48540
rect 60270 48465 60368 48563
rect 60702 48465 60800 48563
rect 61127 48465 61225 48563
rect 12600 48284 12698 48382
rect 54552 48284 54650 48382
rect 6025 48091 6123 48189
rect 6450 48033 6548 48131
rect 6882 48033 6980 48131
rect 7264 48047 7362 48145
rect 7660 48047 7758 48145
rect 12600 48047 12698 48145
rect 54552 48047 54650 48145
rect 59492 48047 59590 48145
rect 59888 48047 59986 48145
rect 60270 48033 60368 48131
rect 60702 48033 60800 48131
rect 61127 48091 61225 48189
rect 12600 47810 12698 47908
rect 54552 47810 54650 47908
rect 6025 47675 6123 47773
rect 6450 47675 6548 47773
rect 6882 47675 6980 47773
rect 7264 47652 7362 47750
rect 7660 47652 7758 47750
rect 59492 47652 59590 47750
rect 59888 47652 59986 47750
rect 60270 47675 60368 47773
rect 60702 47675 60800 47773
rect 61127 47675 61225 47773
rect 12600 47494 12698 47592
rect 54552 47494 54650 47592
rect 6025 47301 6123 47399
rect 6450 47243 6548 47341
rect 6882 47243 6980 47341
rect 7264 47257 7362 47355
rect 7660 47257 7758 47355
rect 12600 47257 12698 47355
rect 54552 47257 54650 47355
rect 59492 47257 59590 47355
rect 59888 47257 59986 47355
rect 60270 47243 60368 47341
rect 60702 47243 60800 47341
rect 61127 47301 61225 47399
rect 12600 47020 12698 47118
rect 54552 47020 54650 47118
rect 6025 46885 6123 46983
rect 6450 46885 6548 46983
rect 6882 46885 6980 46983
rect 7264 46862 7362 46960
rect 7660 46862 7758 46960
rect 59492 46862 59590 46960
rect 59888 46862 59986 46960
rect 60270 46885 60368 46983
rect 60702 46885 60800 46983
rect 61127 46885 61225 46983
rect 12600 46704 12698 46802
rect 54552 46704 54650 46802
rect 6025 46511 6123 46609
rect 6450 46453 6548 46551
rect 6882 46453 6980 46551
rect 7264 46467 7362 46565
rect 7660 46467 7758 46565
rect 12600 46467 12698 46565
rect 54552 46467 54650 46565
rect 59492 46467 59590 46565
rect 59888 46467 59986 46565
rect 60270 46453 60368 46551
rect 60702 46453 60800 46551
rect 61127 46511 61225 46609
rect 12600 46230 12698 46328
rect 54552 46230 54650 46328
rect 6025 46095 6123 46193
rect 6450 46095 6548 46193
rect 6882 46095 6980 46193
rect 7264 46072 7362 46170
rect 7660 46072 7758 46170
rect 59492 46072 59590 46170
rect 59888 46072 59986 46170
rect 60270 46095 60368 46193
rect 60702 46095 60800 46193
rect 61127 46095 61225 46193
rect 12600 45914 12698 46012
rect 54552 45914 54650 46012
rect 6025 45721 6123 45819
rect 6450 45663 6548 45761
rect 6882 45663 6980 45761
rect 7264 45677 7362 45775
rect 7660 45677 7758 45775
rect 12600 45677 12698 45775
rect 54552 45677 54650 45775
rect 59492 45677 59590 45775
rect 59888 45677 59986 45775
rect 60270 45663 60368 45761
rect 60702 45663 60800 45761
rect 61127 45721 61225 45819
rect 12600 45440 12698 45538
rect 54552 45440 54650 45538
rect 6025 45305 6123 45403
rect 6450 45305 6548 45403
rect 6882 45305 6980 45403
rect 7264 45282 7362 45380
rect 7660 45282 7758 45380
rect 59492 45282 59590 45380
rect 59888 45282 59986 45380
rect 60270 45305 60368 45403
rect 60702 45305 60800 45403
rect 61127 45305 61225 45403
rect 12600 45124 12698 45222
rect 54552 45124 54650 45222
rect 6025 44931 6123 45029
rect 6450 44873 6548 44971
rect 6882 44873 6980 44971
rect 7264 44887 7362 44985
rect 7660 44887 7758 44985
rect 12600 44887 12698 44985
rect 54552 44887 54650 44985
rect 59492 44887 59590 44985
rect 59888 44887 59986 44985
rect 60270 44873 60368 44971
rect 60702 44873 60800 44971
rect 61127 44931 61225 45029
rect 12600 44650 12698 44748
rect 54552 44650 54650 44748
rect 6025 44515 6123 44613
rect 6450 44515 6548 44613
rect 6882 44515 6980 44613
rect 7264 44492 7362 44590
rect 7660 44492 7758 44590
rect 59492 44492 59590 44590
rect 59888 44492 59986 44590
rect 60270 44515 60368 44613
rect 60702 44515 60800 44613
rect 61127 44515 61225 44613
rect 12600 44334 12698 44432
rect 54552 44334 54650 44432
rect 6025 44141 6123 44239
rect 6450 44083 6548 44181
rect 6882 44083 6980 44181
rect 7264 44097 7362 44195
rect 7660 44097 7758 44195
rect 12600 44097 12698 44195
rect 54552 44097 54650 44195
rect 59492 44097 59590 44195
rect 59888 44097 59986 44195
rect 60270 44083 60368 44181
rect 60702 44083 60800 44181
rect 61127 44141 61225 44239
rect 12600 43860 12698 43958
rect 54552 43860 54650 43958
rect 6025 43725 6123 43823
rect 6450 43725 6548 43823
rect 6882 43725 6980 43823
rect 7264 43702 7362 43800
rect 7660 43702 7758 43800
rect 59492 43702 59590 43800
rect 59888 43702 59986 43800
rect 60270 43725 60368 43823
rect 60702 43725 60800 43823
rect 61127 43725 61225 43823
rect 12600 43544 12698 43642
rect 54552 43544 54650 43642
rect 6025 43351 6123 43449
rect 6450 43293 6548 43391
rect 6882 43293 6980 43391
rect 7264 43307 7362 43405
rect 7660 43307 7758 43405
rect 12600 43307 12698 43405
rect 54552 43307 54650 43405
rect 59492 43307 59590 43405
rect 59888 43307 59986 43405
rect 60270 43293 60368 43391
rect 60702 43293 60800 43391
rect 61127 43351 61225 43449
rect 12600 43070 12698 43168
rect 54552 43070 54650 43168
rect 6025 42935 6123 43033
rect 6450 42935 6548 43033
rect 6882 42935 6980 43033
rect 7264 42912 7362 43010
rect 7660 42912 7758 43010
rect 59492 42912 59590 43010
rect 59888 42912 59986 43010
rect 60270 42935 60368 43033
rect 60702 42935 60800 43033
rect 61127 42935 61225 43033
rect 12600 42754 12698 42852
rect 54552 42754 54650 42852
rect 6025 42561 6123 42659
rect 6450 42503 6548 42601
rect 6882 42503 6980 42601
rect 7264 42517 7362 42615
rect 7660 42517 7758 42615
rect 12600 42517 12698 42615
rect 54552 42517 54650 42615
rect 59492 42517 59590 42615
rect 59888 42517 59986 42615
rect 60270 42503 60368 42601
rect 60702 42503 60800 42601
rect 61127 42561 61225 42659
rect 12600 42280 12698 42378
rect 54552 42280 54650 42378
rect 6025 42145 6123 42243
rect 6450 42145 6548 42243
rect 6882 42145 6980 42243
rect 7264 42122 7362 42220
rect 7660 42122 7758 42220
rect 59492 42122 59590 42220
rect 59888 42122 59986 42220
rect 60270 42145 60368 42243
rect 60702 42145 60800 42243
rect 61127 42145 61225 42243
rect 12600 41964 12698 42062
rect 54552 41964 54650 42062
rect 6025 41771 6123 41869
rect 6450 41713 6548 41811
rect 6882 41713 6980 41811
rect 7264 41727 7362 41825
rect 7660 41727 7758 41825
rect 12600 41727 12698 41825
rect 54552 41727 54650 41825
rect 59492 41727 59590 41825
rect 59888 41727 59986 41825
rect 60270 41713 60368 41811
rect 60702 41713 60800 41811
rect 61127 41771 61225 41869
rect 12600 41490 12698 41588
rect 54552 41490 54650 41588
rect 6025 41355 6123 41453
rect 6450 41355 6548 41453
rect 6882 41355 6980 41453
rect 7264 41332 7362 41430
rect 7660 41332 7758 41430
rect 59492 41332 59590 41430
rect 59888 41332 59986 41430
rect 60270 41355 60368 41453
rect 60702 41355 60800 41453
rect 61127 41355 61225 41453
rect 12600 41174 12698 41272
rect 54552 41174 54650 41272
rect 6025 40981 6123 41079
rect 6450 40923 6548 41021
rect 6882 40923 6980 41021
rect 7264 40937 7362 41035
rect 7660 40937 7758 41035
rect 12600 40937 12698 41035
rect 54552 40937 54650 41035
rect 59492 40937 59590 41035
rect 59888 40937 59986 41035
rect 60270 40923 60368 41021
rect 60702 40923 60800 41021
rect 61127 40981 61225 41079
rect 12600 40700 12698 40798
rect 54552 40700 54650 40798
rect 6025 40565 6123 40663
rect 6450 40565 6548 40663
rect 6882 40565 6980 40663
rect 7264 40542 7362 40640
rect 7660 40542 7758 40640
rect 59492 40542 59590 40640
rect 59888 40542 59986 40640
rect 60270 40565 60368 40663
rect 60702 40565 60800 40663
rect 61127 40565 61225 40663
rect 12600 40384 12698 40482
rect 54552 40384 54650 40482
rect 6025 40191 6123 40289
rect 6450 40133 6548 40231
rect 6882 40133 6980 40231
rect 7264 40147 7362 40245
rect 7660 40147 7758 40245
rect 12600 40147 12698 40245
rect 54552 40147 54650 40245
rect 59492 40147 59590 40245
rect 59888 40147 59986 40245
rect 60270 40133 60368 40231
rect 60702 40133 60800 40231
rect 61127 40191 61225 40289
rect 12600 39910 12698 40008
rect 54552 39910 54650 40008
rect 6025 39775 6123 39873
rect 6450 39775 6548 39873
rect 6882 39775 6980 39873
rect 7264 39752 7362 39850
rect 7660 39752 7758 39850
rect 59492 39752 59590 39850
rect 59888 39752 59986 39850
rect 60270 39775 60368 39873
rect 60702 39775 60800 39873
rect 61127 39775 61225 39873
rect 12600 39594 12698 39692
rect 54552 39594 54650 39692
rect 6025 39401 6123 39499
rect 6450 39343 6548 39441
rect 6882 39343 6980 39441
rect 7264 39357 7362 39455
rect 7660 39357 7758 39455
rect 12600 39357 12698 39455
rect 54552 39357 54650 39455
rect 59492 39357 59590 39455
rect 59888 39357 59986 39455
rect 60270 39343 60368 39441
rect 60702 39343 60800 39441
rect 61127 39401 61225 39499
rect 12600 39120 12698 39218
rect 54552 39120 54650 39218
rect 6025 38985 6123 39083
rect 6450 38985 6548 39083
rect 6882 38985 6980 39083
rect 7264 38962 7362 39060
rect 7660 38962 7758 39060
rect 59492 38962 59590 39060
rect 59888 38962 59986 39060
rect 60270 38985 60368 39083
rect 60702 38985 60800 39083
rect 61127 38985 61225 39083
rect 12600 38804 12698 38902
rect 54552 38804 54650 38902
rect 6025 38611 6123 38709
rect 6450 38553 6548 38651
rect 6882 38553 6980 38651
rect 7264 38567 7362 38665
rect 7660 38567 7758 38665
rect 12600 38567 12698 38665
rect 54552 38567 54650 38665
rect 59492 38567 59590 38665
rect 59888 38567 59986 38665
rect 60270 38553 60368 38651
rect 60702 38553 60800 38651
rect 61127 38611 61225 38709
rect 12600 38330 12698 38428
rect 54552 38330 54650 38428
rect 6025 38195 6123 38293
rect 6450 38195 6548 38293
rect 6882 38195 6980 38293
rect 7264 38172 7362 38270
rect 7660 38172 7758 38270
rect 59492 38172 59590 38270
rect 59888 38172 59986 38270
rect 60270 38195 60368 38293
rect 60702 38195 60800 38293
rect 61127 38195 61225 38293
rect 12600 38014 12698 38112
rect 54552 38014 54650 38112
rect 6025 37821 6123 37919
rect 6450 37763 6548 37861
rect 6882 37763 6980 37861
rect 7264 37777 7362 37875
rect 7660 37777 7758 37875
rect 12600 37777 12698 37875
rect 54552 37777 54650 37875
rect 59492 37777 59590 37875
rect 59888 37777 59986 37875
rect 60270 37763 60368 37861
rect 60702 37763 60800 37861
rect 61127 37821 61225 37919
rect 12600 37540 12698 37638
rect 54552 37540 54650 37638
rect 6025 37405 6123 37503
rect 6450 37405 6548 37503
rect 6882 37405 6980 37503
rect 7264 37382 7362 37480
rect 7660 37382 7758 37480
rect 59492 37382 59590 37480
rect 59888 37382 59986 37480
rect 60270 37405 60368 37503
rect 60702 37405 60800 37503
rect 61127 37405 61225 37503
rect 12600 37224 12698 37322
rect 54552 37224 54650 37322
rect 6025 37031 6123 37129
rect 6450 36973 6548 37071
rect 6882 36973 6980 37071
rect 7264 36987 7362 37085
rect 7660 36987 7758 37085
rect 12600 36987 12698 37085
rect 54552 36987 54650 37085
rect 59492 36987 59590 37085
rect 59888 36987 59986 37085
rect 60270 36973 60368 37071
rect 60702 36973 60800 37071
rect 61127 37031 61225 37129
rect 12600 36750 12698 36848
rect 54552 36750 54650 36848
rect 6025 36615 6123 36713
rect 6450 36615 6548 36713
rect 6882 36615 6980 36713
rect 7264 36592 7362 36690
rect 7660 36592 7758 36690
rect 59492 36592 59590 36690
rect 59888 36592 59986 36690
rect 60270 36615 60368 36713
rect 60702 36615 60800 36713
rect 61127 36615 61225 36713
rect 12600 36434 12698 36532
rect 54552 36434 54650 36532
rect 6025 36241 6123 36339
rect 6450 36183 6548 36281
rect 6882 36183 6980 36281
rect 7264 36197 7362 36295
rect 7660 36197 7758 36295
rect 12600 36197 12698 36295
rect 54552 36197 54650 36295
rect 59492 36197 59590 36295
rect 59888 36197 59986 36295
rect 60270 36183 60368 36281
rect 60702 36183 60800 36281
rect 61127 36241 61225 36339
rect 12600 35960 12698 36058
rect 54552 35960 54650 36058
rect 6025 35825 6123 35923
rect 6450 35825 6548 35923
rect 6882 35825 6980 35923
rect 7264 35802 7362 35900
rect 7660 35802 7758 35900
rect 59492 35802 59590 35900
rect 59888 35802 59986 35900
rect 60270 35825 60368 35923
rect 60702 35825 60800 35923
rect 61127 35825 61225 35923
rect 12600 35644 12698 35742
rect 54552 35644 54650 35742
rect 6025 35451 6123 35549
rect 6450 35393 6548 35491
rect 6882 35393 6980 35491
rect 7264 35407 7362 35505
rect 7660 35407 7758 35505
rect 8092 35392 8190 35490
rect 8517 35391 8615 35489
rect 9560 35407 9658 35505
rect 11208 35407 11306 35505
rect 12600 35407 12698 35505
rect 54552 35407 54650 35505
rect 55944 35407 56042 35505
rect 57592 35407 57690 35505
rect 58635 35391 58733 35489
rect 59060 35392 59158 35490
rect 59492 35407 59590 35505
rect 59888 35407 59986 35505
rect 60270 35393 60368 35491
rect 60702 35393 60800 35491
rect 61127 35451 61225 35549
rect 12600 35170 12698 35268
rect 54552 35170 54650 35268
rect 6025 35035 6123 35133
rect 6450 35035 6548 35133
rect 6882 35035 6980 35133
rect 7264 35012 7362 35110
rect 7660 35012 7758 35110
rect 59492 35012 59590 35110
rect 59888 35012 59986 35110
rect 60270 35035 60368 35133
rect 60702 35035 60800 35133
rect 61127 35035 61225 35133
rect 12600 34854 12698 34952
rect 54552 34854 54650 34952
rect 6025 34661 6123 34759
rect 6450 34603 6548 34701
rect 6882 34603 6980 34701
rect 7264 34617 7362 34715
rect 7660 34617 7758 34715
rect 12600 34617 12698 34715
rect 54552 34617 54650 34715
rect 59492 34617 59590 34715
rect 59888 34617 59986 34715
rect 60270 34603 60368 34701
rect 60702 34603 60800 34701
rect 61127 34661 61225 34759
rect 12600 34380 12698 34478
rect 54552 34380 54650 34478
rect 6025 34245 6123 34343
rect 6450 34245 6548 34343
rect 6882 34245 6980 34343
rect 7264 34222 7362 34320
rect 7660 34222 7758 34320
rect 59492 34222 59590 34320
rect 59888 34222 59986 34320
rect 60270 34245 60368 34343
rect 60702 34245 60800 34343
rect 61127 34245 61225 34343
rect 12600 34064 12698 34162
rect 54552 34064 54650 34162
rect 6025 33871 6123 33969
rect 6450 33813 6548 33911
rect 6882 33813 6980 33911
rect 7264 33827 7362 33925
rect 7660 33827 7758 33925
rect 12600 33827 12698 33925
rect 54552 33827 54650 33925
rect 59492 33827 59590 33925
rect 59888 33827 59986 33925
rect 60270 33813 60368 33911
rect 60702 33813 60800 33911
rect 61127 33871 61225 33969
rect 12600 33590 12698 33688
rect 54552 33590 54650 33688
rect 6025 33455 6123 33553
rect 6450 33455 6548 33553
rect 6882 33455 6980 33553
rect 7264 33432 7362 33530
rect 7660 33432 7758 33530
rect 59492 33432 59590 33530
rect 59888 33432 59986 33530
rect 60270 33455 60368 33553
rect 60702 33455 60800 33553
rect 61127 33455 61225 33553
rect 12600 33274 12698 33372
rect 54552 33274 54650 33372
rect 6025 33081 6123 33179
rect 6450 33023 6548 33121
rect 6882 33023 6980 33121
rect 7264 33037 7362 33135
rect 7660 33037 7758 33135
rect 12600 33037 12698 33135
rect 54552 33037 54650 33135
rect 59492 33037 59590 33135
rect 59888 33037 59986 33135
rect 60270 33023 60368 33121
rect 60702 33023 60800 33121
rect 61127 33081 61225 33179
rect 12600 32800 12698 32898
rect 54552 32800 54650 32898
rect 6025 32665 6123 32763
rect 6450 32665 6548 32763
rect 6882 32665 6980 32763
rect 7264 32642 7362 32740
rect 7660 32642 7758 32740
rect 59492 32642 59590 32740
rect 59888 32642 59986 32740
rect 60270 32665 60368 32763
rect 60702 32665 60800 32763
rect 61127 32665 61225 32763
rect 12600 32484 12698 32582
rect 54552 32484 54650 32582
rect 6025 32291 6123 32389
rect 6450 32233 6548 32331
rect 6882 32233 6980 32331
rect 7264 32247 7362 32345
rect 7660 32247 7758 32345
rect 12600 32247 12698 32345
rect 54552 32247 54650 32345
rect 59492 32247 59590 32345
rect 59888 32247 59986 32345
rect 60270 32233 60368 32331
rect 60702 32233 60800 32331
rect 61127 32291 61225 32389
rect 12600 32010 12698 32108
rect 54552 32010 54650 32108
rect 6025 31875 6123 31973
rect 6450 31875 6548 31973
rect 6882 31875 6980 31973
rect 7264 31852 7362 31950
rect 7660 31852 7758 31950
rect 59492 31852 59590 31950
rect 59888 31852 59986 31950
rect 60270 31875 60368 31973
rect 60702 31875 60800 31973
rect 61127 31875 61225 31973
rect 12600 31694 12698 31792
rect 54552 31694 54650 31792
rect 6025 31501 6123 31599
rect 6450 31443 6548 31541
rect 6882 31443 6980 31541
rect 7264 31457 7362 31555
rect 7660 31457 7758 31555
rect 12600 31457 12698 31555
rect 54552 31457 54650 31555
rect 59492 31457 59590 31555
rect 59888 31457 59986 31555
rect 60270 31443 60368 31541
rect 60702 31443 60800 31541
rect 61127 31501 61225 31599
rect 12600 31220 12698 31318
rect 54552 31220 54650 31318
rect 6025 31085 6123 31183
rect 6450 31085 6548 31183
rect 6882 31085 6980 31183
rect 7264 31062 7362 31160
rect 7660 31062 7758 31160
rect 59492 31062 59590 31160
rect 59888 31062 59986 31160
rect 60270 31085 60368 31183
rect 60702 31085 60800 31183
rect 61127 31085 61225 31183
rect 12600 30904 12698 31002
rect 54552 30904 54650 31002
rect 6025 30711 6123 30809
rect 6450 30653 6548 30751
rect 6882 30653 6980 30751
rect 7264 30667 7362 30765
rect 7660 30667 7758 30765
rect 12600 30667 12698 30765
rect 54552 30667 54650 30765
rect 59492 30667 59590 30765
rect 59888 30667 59986 30765
rect 60270 30653 60368 30751
rect 60702 30653 60800 30751
rect 61127 30711 61225 30809
rect 12600 30430 12698 30528
rect 54552 30430 54650 30528
rect 6025 30295 6123 30393
rect 6450 30295 6548 30393
rect 6882 30295 6980 30393
rect 7264 30272 7362 30370
rect 7660 30272 7758 30370
rect 59492 30272 59590 30370
rect 59888 30272 59986 30370
rect 60270 30295 60368 30393
rect 60702 30295 60800 30393
rect 61127 30295 61225 30393
rect 12600 30114 12698 30212
rect 54552 30114 54650 30212
rect 6025 29921 6123 30019
rect 6450 29863 6548 29961
rect 6882 29863 6980 29961
rect 7264 29877 7362 29975
rect 7660 29877 7758 29975
rect 12600 29877 12698 29975
rect 54552 29877 54650 29975
rect 59492 29877 59590 29975
rect 59888 29877 59986 29975
rect 60270 29863 60368 29961
rect 60702 29863 60800 29961
rect 61127 29921 61225 30019
rect 12600 29640 12698 29738
rect 54552 29640 54650 29738
rect 6025 29505 6123 29603
rect 6450 29505 6548 29603
rect 6882 29505 6980 29603
rect 7264 29482 7362 29580
rect 7660 29482 7758 29580
rect 59492 29482 59590 29580
rect 59888 29482 59986 29580
rect 60270 29505 60368 29603
rect 60702 29505 60800 29603
rect 61127 29505 61225 29603
rect 12600 29324 12698 29422
rect 54552 29324 54650 29422
rect 6025 29131 6123 29229
rect 6450 29073 6548 29171
rect 6882 29073 6980 29171
rect 7264 29087 7362 29185
rect 7660 29087 7758 29185
rect 12600 29087 12698 29185
rect 54552 29087 54650 29185
rect 59492 29087 59590 29185
rect 59888 29087 59986 29185
rect 60270 29073 60368 29171
rect 60702 29073 60800 29171
rect 61127 29131 61225 29229
rect 12600 28850 12698 28948
rect 54552 28850 54650 28948
rect 6025 28715 6123 28813
rect 6450 28715 6548 28813
rect 6882 28715 6980 28813
rect 7264 28692 7362 28790
rect 7660 28692 7758 28790
rect 59492 28692 59590 28790
rect 59888 28692 59986 28790
rect 60270 28715 60368 28813
rect 60702 28715 60800 28813
rect 61127 28715 61225 28813
rect 12600 28534 12698 28632
rect 54552 28534 54650 28632
rect 6025 28341 6123 28439
rect 6450 28283 6548 28381
rect 6882 28283 6980 28381
rect 7264 28297 7362 28395
rect 7660 28297 7758 28395
rect 12600 28297 12698 28395
rect 54552 28297 54650 28395
rect 59492 28297 59590 28395
rect 59888 28297 59986 28395
rect 60270 28283 60368 28381
rect 60702 28283 60800 28381
rect 61127 28341 61225 28439
rect 12600 28060 12698 28158
rect 54552 28060 54650 28158
rect 6025 27925 6123 28023
rect 6450 27925 6548 28023
rect 6882 27925 6980 28023
rect 7264 27902 7362 28000
rect 7660 27902 7758 28000
rect 59492 27902 59590 28000
rect 59888 27902 59986 28000
rect 60270 27925 60368 28023
rect 60702 27925 60800 28023
rect 61127 27925 61225 28023
rect 12600 27744 12698 27842
rect 54552 27744 54650 27842
rect 6025 27551 6123 27649
rect 6450 27493 6548 27591
rect 6882 27493 6980 27591
rect 7264 27507 7362 27605
rect 7660 27507 7758 27605
rect 12600 27507 12698 27605
rect 54552 27507 54650 27605
rect 59492 27507 59590 27605
rect 59888 27507 59986 27605
rect 60270 27493 60368 27591
rect 60702 27493 60800 27591
rect 61127 27551 61225 27649
rect 12600 27270 12698 27368
rect 54552 27270 54650 27368
rect 6025 27135 6123 27233
rect 6450 27135 6548 27233
rect 6882 27135 6980 27233
rect 7264 27112 7362 27210
rect 7660 27112 7758 27210
rect 59492 27112 59590 27210
rect 59888 27112 59986 27210
rect 60270 27135 60368 27233
rect 60702 27135 60800 27233
rect 61127 27135 61225 27233
rect 12600 26954 12698 27052
rect 54552 26954 54650 27052
rect 6025 26761 6123 26859
rect 6450 26703 6548 26801
rect 6882 26703 6980 26801
rect 7264 26717 7362 26815
rect 7660 26717 7758 26815
rect 12600 26717 12698 26815
rect 54552 26717 54650 26815
rect 59492 26717 59590 26815
rect 59888 26717 59986 26815
rect 60270 26703 60368 26801
rect 60702 26703 60800 26801
rect 61127 26761 61225 26859
rect 12600 26480 12698 26578
rect 54552 26480 54650 26578
rect 6025 26345 6123 26443
rect 6450 26345 6548 26443
rect 6882 26345 6980 26443
rect 7264 26322 7362 26420
rect 7660 26322 7758 26420
rect 59492 26322 59590 26420
rect 59888 26322 59986 26420
rect 60270 26345 60368 26443
rect 60702 26345 60800 26443
rect 61127 26345 61225 26443
rect 12600 26164 12698 26262
rect 54552 26164 54650 26262
rect 6025 25971 6123 26069
rect 6450 25913 6548 26011
rect 6882 25913 6980 26011
rect 7264 25927 7362 26025
rect 7660 25927 7758 26025
rect 12600 25927 12698 26025
rect 54552 25927 54650 26025
rect 59492 25927 59590 26025
rect 59888 25927 59986 26025
rect 60270 25913 60368 26011
rect 60702 25913 60800 26011
rect 61127 25971 61225 26069
rect 12600 25690 12698 25788
rect 54552 25690 54650 25788
rect 6025 25555 6123 25653
rect 6450 25555 6548 25653
rect 6882 25555 6980 25653
rect 7264 25532 7362 25630
rect 7660 25532 7758 25630
rect 59492 25532 59590 25630
rect 59888 25532 59986 25630
rect 60270 25555 60368 25653
rect 60702 25555 60800 25653
rect 61127 25555 61225 25653
rect 12600 25374 12698 25472
rect 54552 25374 54650 25472
rect 6025 25181 6123 25279
rect 6450 25123 6548 25221
rect 6882 25123 6980 25221
rect 7264 25137 7362 25235
rect 7660 25137 7758 25235
rect 12600 25137 12698 25235
rect 54552 25137 54650 25235
rect 59492 25137 59590 25235
rect 59888 25137 59986 25235
rect 60270 25123 60368 25221
rect 60702 25123 60800 25221
rect 61127 25181 61225 25279
rect 12600 24900 12698 24998
rect 54552 24900 54650 24998
rect 6025 24765 6123 24863
rect 6450 24765 6548 24863
rect 6882 24765 6980 24863
rect 7264 24742 7362 24840
rect 7660 24742 7758 24840
rect 59492 24742 59590 24840
rect 59888 24742 59986 24840
rect 60270 24765 60368 24863
rect 60702 24765 60800 24863
rect 61127 24765 61225 24863
rect 12600 24584 12698 24682
rect 54552 24584 54650 24682
rect 6025 24391 6123 24489
rect 6450 24333 6548 24431
rect 6882 24333 6980 24431
rect 7264 24347 7362 24445
rect 7660 24347 7758 24445
rect 12600 24347 12698 24445
rect 54552 24347 54650 24445
rect 59492 24347 59590 24445
rect 59888 24347 59986 24445
rect 60270 24333 60368 24431
rect 60702 24333 60800 24431
rect 61127 24391 61225 24489
rect 12600 24110 12698 24208
rect 54552 24110 54650 24208
rect 6025 23975 6123 24073
rect 6450 23975 6548 24073
rect 6882 23975 6980 24073
rect 7264 23952 7362 24050
rect 7660 23952 7758 24050
rect 59492 23952 59590 24050
rect 59888 23952 59986 24050
rect 60270 23975 60368 24073
rect 60702 23975 60800 24073
rect 61127 23975 61225 24073
rect 12600 23794 12698 23892
rect 54552 23794 54650 23892
rect 6025 23601 6123 23699
rect 6450 23543 6548 23641
rect 6882 23543 6980 23641
rect 7264 23557 7362 23655
rect 7660 23557 7758 23655
rect 12600 23557 12698 23655
rect 54552 23557 54650 23655
rect 59492 23557 59590 23655
rect 59888 23557 59986 23655
rect 60270 23543 60368 23641
rect 60702 23543 60800 23641
rect 61127 23601 61225 23699
rect 12600 23320 12698 23418
rect 54552 23320 54650 23418
rect 6025 23185 6123 23283
rect 6450 23185 6548 23283
rect 6882 23185 6980 23283
rect 7264 23162 7362 23260
rect 7660 23162 7758 23260
rect 59492 23162 59590 23260
rect 59888 23162 59986 23260
rect 60270 23185 60368 23283
rect 60702 23185 60800 23283
rect 61127 23185 61225 23283
rect 12600 23004 12698 23102
rect 54552 23004 54650 23102
rect 6025 22811 6123 22909
rect 6450 22753 6548 22851
rect 6882 22753 6980 22851
rect 7264 22767 7362 22865
rect 7660 22767 7758 22865
rect 12600 22767 12698 22865
rect 54552 22767 54650 22865
rect 59492 22767 59590 22865
rect 59888 22767 59986 22865
rect 60270 22753 60368 22851
rect 60702 22753 60800 22851
rect 61127 22811 61225 22909
rect 12600 22530 12698 22628
rect 54552 22530 54650 22628
rect 6025 22395 6123 22493
rect 6450 22395 6548 22493
rect 6882 22395 6980 22493
rect 7264 22372 7362 22470
rect 7660 22372 7758 22470
rect 59492 22372 59590 22470
rect 59888 22372 59986 22470
rect 60270 22395 60368 22493
rect 60702 22395 60800 22493
rect 61127 22395 61225 22493
rect 12600 22214 12698 22312
rect 54552 22214 54650 22312
rect 6025 22021 6123 22119
rect 6450 21963 6548 22061
rect 6882 21963 6980 22061
rect 7264 21977 7362 22075
rect 7660 21977 7758 22075
rect 12600 21977 12698 22075
rect 54552 21977 54650 22075
rect 59492 21977 59590 22075
rect 59888 21977 59986 22075
rect 60270 21963 60368 22061
rect 60702 21963 60800 22061
rect 61127 22021 61225 22119
rect 12600 21740 12698 21838
rect 54552 21740 54650 21838
rect 6025 21605 6123 21703
rect 6450 21605 6548 21703
rect 6882 21605 6980 21703
rect 7264 21582 7362 21680
rect 7660 21582 7758 21680
rect 59492 21582 59590 21680
rect 59888 21582 59986 21680
rect 60270 21605 60368 21703
rect 60702 21605 60800 21703
rect 61127 21605 61225 21703
rect 12600 21424 12698 21522
rect 54552 21424 54650 21522
rect 6025 21231 6123 21329
rect 6450 21173 6548 21271
rect 6882 21173 6980 21271
rect 7264 21187 7362 21285
rect 7660 21187 7758 21285
rect 12600 21187 12698 21285
rect 54552 21187 54650 21285
rect 59492 21187 59590 21285
rect 59888 21187 59986 21285
rect 60270 21173 60368 21271
rect 60702 21173 60800 21271
rect 61127 21231 61225 21329
rect 12600 20950 12698 21048
rect 54552 20950 54650 21048
rect 6025 20815 6123 20913
rect 6450 20815 6548 20913
rect 6882 20815 6980 20913
rect 7264 20792 7362 20890
rect 7660 20792 7758 20890
rect 59492 20792 59590 20890
rect 59888 20792 59986 20890
rect 60270 20815 60368 20913
rect 60702 20815 60800 20913
rect 61127 20815 61225 20913
rect 12600 20634 12698 20732
rect 54552 20634 54650 20732
rect 6025 20441 6123 20539
rect 6450 20383 6548 20481
rect 6882 20383 6980 20481
rect 7264 20397 7362 20495
rect 7660 20397 7758 20495
rect 12600 20397 12698 20495
rect 54552 20397 54650 20495
rect 59492 20397 59590 20495
rect 59888 20397 59986 20495
rect 60270 20383 60368 20481
rect 60702 20383 60800 20481
rect 61127 20441 61225 20539
rect 12600 20160 12698 20258
rect 54552 20160 54650 20258
rect 6025 20025 6123 20123
rect 6450 20025 6548 20123
rect 6882 20025 6980 20123
rect 7264 20002 7362 20100
rect 7660 20002 7758 20100
rect 59492 20002 59590 20100
rect 59888 20002 59986 20100
rect 60270 20025 60368 20123
rect 60702 20025 60800 20123
rect 61127 20025 61225 20123
rect 12600 19844 12698 19942
rect 54552 19844 54650 19942
rect 6025 19651 6123 19749
rect 6450 19593 6548 19691
rect 6882 19593 6980 19691
rect 7264 19607 7362 19705
rect 7660 19607 7758 19705
rect 12600 19607 12698 19705
rect 54552 19607 54650 19705
rect 59492 19607 59590 19705
rect 59888 19607 59986 19705
rect 60270 19593 60368 19691
rect 60702 19593 60800 19691
rect 61127 19651 61225 19749
rect 12600 19370 12698 19468
rect 54552 19370 54650 19468
rect 6025 19235 6123 19333
rect 6450 19235 6548 19333
rect 6882 19235 6980 19333
rect 7264 19212 7362 19310
rect 7660 19212 7758 19310
rect 59492 19212 59590 19310
rect 59888 19212 59986 19310
rect 60270 19235 60368 19333
rect 60702 19235 60800 19333
rect 61127 19235 61225 19333
rect 12600 19054 12698 19152
rect 54552 19054 54650 19152
rect 6025 18861 6123 18959
rect 6450 18803 6548 18901
rect 6882 18803 6980 18901
rect 7264 18817 7362 18915
rect 7660 18817 7758 18915
rect 12600 18817 12698 18915
rect 54552 18817 54650 18915
rect 59492 18817 59590 18915
rect 59888 18817 59986 18915
rect 60270 18803 60368 18901
rect 60702 18803 60800 18901
rect 61127 18861 61225 18959
rect 12600 18580 12698 18678
rect 54552 18580 54650 18678
rect 6025 18445 6123 18543
rect 6450 18445 6548 18543
rect 6882 18445 6980 18543
rect 7264 18422 7362 18520
rect 7660 18422 7758 18520
rect 59492 18422 59590 18520
rect 59888 18422 59986 18520
rect 60270 18445 60368 18543
rect 60702 18445 60800 18543
rect 61127 18445 61225 18543
rect 12600 18264 12698 18362
rect 54552 18264 54650 18362
rect 6025 18071 6123 18169
rect 6450 18013 6548 18111
rect 6882 18013 6980 18111
rect 7264 18027 7362 18125
rect 7660 18027 7758 18125
rect 12600 18027 12698 18125
rect 54552 18027 54650 18125
rect 59492 18027 59590 18125
rect 59888 18027 59986 18125
rect 60270 18013 60368 18111
rect 60702 18013 60800 18111
rect 61127 18071 61225 18169
rect 12600 17790 12698 17888
rect 54552 17790 54650 17888
rect 2611 17655 2709 17753
rect 3036 17655 3134 17753
rect 3468 17655 3566 17753
rect 3850 17632 3948 17730
rect 4246 17632 4344 17730
rect 6025 17655 6123 17753
rect 6450 17655 6548 17753
rect 6882 17655 6980 17753
rect 7264 17632 7362 17730
rect 7660 17632 7758 17730
rect 59492 17632 59590 17730
rect 59888 17632 59986 17730
rect 60270 17655 60368 17753
rect 60702 17655 60800 17753
rect 61127 17655 61225 17753
rect 62906 17632 63004 17730
rect 63302 17632 63400 17730
rect 63684 17655 63782 17753
rect 64116 17655 64214 17753
rect 64541 17655 64639 17753
rect 12600 17474 12698 17572
rect 54552 17474 54650 17572
rect 6025 17281 6123 17379
rect 6450 17223 6548 17321
rect 6882 17223 6980 17321
rect 7264 17237 7362 17335
rect 7660 17237 7758 17335
rect 12600 17237 12698 17335
rect 54552 17237 54650 17335
rect 59492 17237 59590 17335
rect 59888 17237 59986 17335
rect 60270 17223 60368 17321
rect 60702 17223 60800 17321
rect 61127 17281 61225 17379
rect 12600 17000 12698 17098
rect 54552 17000 54650 17098
rect 2611 16865 2709 16963
rect 3036 16865 3134 16963
rect 3468 16865 3566 16963
rect 3850 16842 3948 16940
rect 4246 16842 4344 16940
rect 6025 16865 6123 16963
rect 6450 16865 6548 16963
rect 6882 16865 6980 16963
rect 7264 16842 7362 16940
rect 7660 16842 7758 16940
rect 59492 16842 59590 16940
rect 59888 16842 59986 16940
rect 60270 16865 60368 16963
rect 60702 16865 60800 16963
rect 61127 16865 61225 16963
rect 62906 16842 63004 16940
rect 63302 16842 63400 16940
rect 63684 16865 63782 16963
rect 64116 16865 64214 16963
rect 64541 16865 64639 16963
rect 12600 16684 12698 16782
rect 54552 16684 54650 16782
rect 6025 16491 6123 16589
rect 6450 16433 6548 16531
rect 6882 16433 6980 16531
rect 7264 16447 7362 16545
rect 7660 16447 7758 16545
rect 12600 16447 12698 16545
rect 54552 16447 54650 16545
rect 59492 16447 59590 16545
rect 59888 16447 59986 16545
rect 60270 16433 60368 16531
rect 60702 16433 60800 16531
rect 61127 16491 61225 16589
rect 12600 16210 12698 16308
rect 54552 16210 54650 16308
rect 2611 16075 2709 16173
rect 3036 16075 3134 16173
rect 3468 16075 3566 16173
rect 3850 16052 3948 16150
rect 4246 16052 4344 16150
rect 6025 16075 6123 16173
rect 6450 16075 6548 16173
rect 6882 16075 6980 16173
rect 7264 16052 7362 16150
rect 7660 16052 7758 16150
rect 59492 16052 59590 16150
rect 59888 16052 59986 16150
rect 60270 16075 60368 16173
rect 60702 16075 60800 16173
rect 61127 16075 61225 16173
rect 62906 16052 63004 16150
rect 63302 16052 63400 16150
rect 63684 16075 63782 16173
rect 64116 16075 64214 16173
rect 64541 16075 64639 16173
rect 12600 15894 12698 15992
rect 54552 15894 54650 15992
rect 6025 15701 6123 15799
rect 6450 15643 6548 15741
rect 6882 15643 6980 15741
rect 7264 15657 7362 15755
rect 7660 15657 7758 15755
rect 12600 15657 12698 15755
rect 54552 15657 54650 15755
rect 59492 15657 59590 15755
rect 59888 15657 59986 15755
rect 60270 15643 60368 15741
rect 60702 15643 60800 15741
rect 61127 15701 61225 15799
rect 12600 15420 12698 15518
rect 54552 15420 54650 15518
rect 1156 15262 1254 15360
rect 1552 15262 1650 15360
rect 2611 15285 2709 15383
rect 3036 15285 3134 15383
rect 3468 15285 3566 15383
rect 3850 15262 3948 15360
rect 4246 15262 4344 15360
rect 6025 15285 6123 15383
rect 6450 15285 6548 15383
rect 6882 15285 6980 15383
rect 7264 15262 7362 15360
rect 7660 15262 7758 15360
rect 59492 15262 59590 15360
rect 59888 15262 59986 15360
rect 60270 15285 60368 15383
rect 60702 15285 60800 15383
rect 61127 15285 61225 15383
rect 62906 15262 63004 15360
rect 63302 15262 63400 15360
rect 63684 15285 63782 15383
rect 64116 15285 64214 15383
rect 64541 15285 64639 15383
rect 65600 15262 65698 15360
rect 65996 15262 66094 15360
rect 12600 15104 12698 15202
rect 54552 15104 54650 15202
rect 6025 14911 6123 15009
rect 6450 14853 6548 14951
rect 6882 14853 6980 14951
rect 7264 14867 7362 14965
rect 7660 14867 7758 14965
rect 12600 14867 12698 14965
rect 54552 14867 54650 14965
rect 59492 14867 59590 14965
rect 59888 14867 59986 14965
rect 60270 14853 60368 14951
rect 60702 14853 60800 14951
rect 61127 14911 61225 15009
rect 12600 14630 12698 14728
rect 54552 14630 54650 14728
rect 6025 14495 6123 14593
rect 6450 14495 6548 14593
rect 6882 14495 6980 14593
rect 7264 14472 7362 14570
rect 7660 14472 7758 14570
rect 59492 14472 59590 14570
rect 59888 14472 59986 14570
rect 60270 14495 60368 14593
rect 60702 14495 60800 14593
rect 61127 14495 61225 14593
rect 12600 14314 12698 14412
rect 54552 14314 54650 14412
rect 6025 14121 6123 14219
rect 6450 14063 6548 14161
rect 6882 14063 6980 14161
rect 7264 14077 7362 14175
rect 7660 14077 7758 14175
rect 12600 14077 12698 14175
rect 54552 14077 54650 14175
rect 59492 14077 59590 14175
rect 59888 14077 59986 14175
rect 60270 14063 60368 14161
rect 60702 14063 60800 14161
rect 61127 14121 61225 14219
rect 12600 13840 12698 13938
rect 54552 13840 54650 13938
rect 3046 13689 3144 13787
rect 3471 13689 3569 13787
rect 3850 13682 3948 13780
rect 4246 13682 4344 13780
rect 6025 13705 6123 13803
rect 6450 13705 6548 13803
rect 6882 13705 6980 13803
rect 7264 13682 7362 13780
rect 7660 13682 7758 13780
rect 59492 13682 59590 13780
rect 59888 13682 59986 13780
rect 60270 13705 60368 13803
rect 60702 13705 60800 13803
rect 61127 13705 61225 13803
rect 62906 13682 63004 13780
rect 63302 13682 63400 13780
rect 63681 13689 63779 13787
rect 64106 13689 64204 13787
rect 12600 13524 12698 13622
rect 54552 13524 54650 13622
rect 6025 13331 6123 13429
rect 6450 13273 6548 13371
rect 6882 13273 6980 13371
rect 7264 13287 7362 13385
rect 7660 13287 7758 13385
rect 12600 13287 12698 13385
rect 54552 13287 54650 13385
rect 59492 13287 59590 13385
rect 59888 13287 59986 13385
rect 60270 13273 60368 13371
rect 60702 13273 60800 13371
rect 61127 13331 61225 13429
rect 12600 13050 12698 13148
rect 54552 13050 54650 13148
rect 1752 12892 1850 12990
rect 2148 12892 2246 12990
rect 3046 12899 3144 12997
rect 3471 12899 3569 12997
rect 3850 12892 3948 12990
rect 4246 12892 4344 12990
rect 6025 12915 6123 13013
rect 6450 12915 6548 13013
rect 6882 12915 6980 13013
rect 7264 12892 7362 12990
rect 7660 12892 7758 12990
rect 59492 12892 59590 12990
rect 59888 12892 59986 12990
rect 60270 12915 60368 13013
rect 60702 12915 60800 13013
rect 61127 12915 61225 13013
rect 62906 12892 63004 12990
rect 63302 12892 63400 12990
rect 63681 12899 63779 12997
rect 64106 12899 64204 12997
rect 65004 12892 65102 12990
rect 65400 12892 65498 12990
rect 12600 12734 12698 12832
rect 54552 12734 54650 12832
rect 6025 12541 6123 12639
rect 6450 12483 6548 12581
rect 6882 12483 6980 12581
rect 7264 12497 7362 12595
rect 7660 12497 7758 12595
rect 12600 12497 12698 12595
rect 54552 12497 54650 12595
rect 59492 12497 59590 12595
rect 59888 12497 59986 12595
rect 60270 12483 60368 12581
rect 60702 12483 60800 12581
rect 61127 12541 61225 12639
rect 12600 12260 12698 12358
rect 54552 12260 54650 12358
rect 6025 12125 6123 12223
rect 6450 12125 6548 12223
rect 6882 12125 6980 12223
rect 7264 12102 7362 12200
rect 7660 12102 7758 12200
rect 59492 12102 59590 12200
rect 59888 12102 59986 12200
rect 60270 12125 60368 12223
rect 60702 12125 60800 12223
rect 61127 12125 61225 12223
rect 12600 11944 12698 12042
rect 54552 11944 54650 12042
rect 6025 11751 6123 11849
rect 6450 11693 6548 11791
rect 6882 11693 6980 11791
rect 7264 11707 7362 11805
rect 7660 11707 7758 11805
rect 12600 11707 12698 11805
rect 54552 11707 54650 11805
rect 59492 11707 59590 11805
rect 59888 11707 59986 11805
rect 60270 11693 60368 11791
rect 60702 11693 60800 11791
rect 61127 11751 61225 11849
rect 12600 11470 12698 11568
rect 54552 11470 54650 11568
rect 3046 11319 3144 11417
rect 3471 11319 3569 11417
rect 3850 11312 3948 11410
rect 4246 11312 4344 11410
rect 6025 11335 6123 11433
rect 6450 11335 6548 11433
rect 6882 11335 6980 11433
rect 7264 11312 7362 11410
rect 7660 11312 7758 11410
rect 59492 11312 59590 11410
rect 59888 11312 59986 11410
rect 60270 11335 60368 11433
rect 60702 11335 60800 11433
rect 61127 11335 61225 11433
rect 62906 11312 63004 11410
rect 63302 11312 63400 11410
rect 63681 11319 63779 11417
rect 64106 11319 64204 11417
rect 12600 11154 12698 11252
rect 54552 11154 54650 11252
rect 6025 10961 6123 11059
rect 6450 10903 6548 11001
rect 6882 10903 6980 11001
rect 7264 10917 7362 11015
rect 7660 10917 7758 11015
rect 12600 10917 12698 11015
rect 54552 10917 54650 11015
rect 59492 10917 59590 11015
rect 59888 10917 59986 11015
rect 60270 10903 60368 11001
rect 60702 10903 60800 11001
rect 61127 10961 61225 11059
rect 12600 10680 12698 10778
rect 54552 10680 54650 10778
rect 1752 10522 1850 10620
rect 2148 10522 2246 10620
rect 3046 10529 3144 10627
rect 3471 10529 3569 10627
rect 3850 10522 3948 10620
rect 4246 10522 4344 10620
rect 6025 10545 6123 10643
rect 6450 10545 6548 10643
rect 6882 10545 6980 10643
rect 7264 10522 7362 10620
rect 7660 10522 7758 10620
rect 59492 10522 59590 10620
rect 59888 10522 59986 10620
rect 60270 10545 60368 10643
rect 60702 10545 60800 10643
rect 61127 10545 61225 10643
rect 62906 10522 63004 10620
rect 63302 10522 63400 10620
rect 63681 10529 63779 10627
rect 64106 10529 64204 10627
rect 65004 10522 65102 10620
rect 65400 10522 65498 10620
rect 12600 10364 12698 10462
rect 54552 10364 54650 10462
rect 12600 10127 12698 10225
rect 54552 10127 54650 10225
rect 7685 9936 7783 10034
rect 8517 9942 8615 10040
rect 11208 9930 11306 10028
rect 12234 10000 12332 10098
rect 54918 10000 55016 10098
rect 13296 9566 13394 9664
rect 13920 9566 14018 9664
rect 14544 9566 14642 9664
rect 15168 9566 15266 9664
rect 15792 9566 15890 9664
rect 16416 9566 16514 9664
rect 17040 9566 17138 9664
rect 17664 9566 17762 9664
rect 18288 9566 18386 9664
rect 18912 9566 19010 9664
rect 19536 9566 19634 9664
rect 20160 9566 20258 9664
rect 20784 9566 20882 9664
rect 21408 9566 21506 9664
rect 22032 9566 22130 9664
rect 22656 9566 22754 9664
rect 23280 9566 23378 9664
rect 23904 9566 24002 9664
rect 24528 9566 24626 9664
rect 25152 9566 25250 9664
rect 25776 9566 25874 9664
rect 26400 9566 26498 9664
rect 27024 9566 27122 9664
rect 27648 9566 27746 9664
rect 28272 9566 28370 9664
rect 28896 9566 28994 9664
rect 29520 9566 29618 9664
rect 30144 9566 30242 9664
rect 30768 9566 30866 9664
rect 31392 9566 31490 9664
rect 32016 9566 32114 9664
rect 32640 9566 32738 9664
rect 33264 9566 33362 9664
rect 33888 9566 33986 9664
rect 34512 9566 34610 9664
rect 35136 9566 35234 9664
rect 35760 9566 35858 9664
rect 36384 9566 36482 9664
rect 37008 9566 37106 9664
rect 37632 9566 37730 9664
rect 38256 9566 38354 9664
rect 38880 9566 38978 9664
rect 39504 9566 39602 9664
rect 40128 9566 40226 9664
rect 40752 9566 40850 9664
rect 41376 9566 41474 9664
rect 42000 9566 42098 9664
rect 42624 9566 42722 9664
rect 43248 9566 43346 9664
rect 43872 9566 43970 9664
rect 44496 9566 44594 9664
rect 45120 9566 45218 9664
rect 45744 9566 45842 9664
rect 46368 9566 46466 9664
rect 46992 9566 47090 9664
rect 47616 9566 47714 9664
rect 48240 9566 48338 9664
rect 48864 9566 48962 9664
rect 49488 9566 49586 9664
rect 50112 9566 50210 9664
rect 50736 9566 50834 9664
rect 51360 9566 51458 9664
rect 51984 9566 52082 9664
rect 52608 9566 52706 9664
rect 53232 9566 53330 9664
rect 53856 9566 53954 9664
rect 13415 8975 13513 9073
rect 13801 8975 13899 9073
rect 14663 8975 14761 9073
rect 15049 8975 15147 9073
rect 15911 8975 16009 9073
rect 16297 8975 16395 9073
rect 17159 8975 17257 9073
rect 17545 8975 17643 9073
rect 18407 8975 18505 9073
rect 18793 8975 18891 9073
rect 19655 8975 19753 9073
rect 20041 8975 20139 9073
rect 20903 8975 21001 9073
rect 21289 8975 21387 9073
rect 22151 8975 22249 9073
rect 22537 8975 22635 9073
rect 23399 8975 23497 9073
rect 23785 8975 23883 9073
rect 24647 8975 24745 9073
rect 25033 8975 25131 9073
rect 25895 8975 25993 9073
rect 26281 8975 26379 9073
rect 27143 8975 27241 9073
rect 27529 8975 27627 9073
rect 28391 8975 28489 9073
rect 28777 8975 28875 9073
rect 29639 8975 29737 9073
rect 30025 8975 30123 9073
rect 30887 8975 30985 9073
rect 31273 8975 31371 9073
rect 32135 8975 32233 9073
rect 32521 8975 32619 9073
rect 33383 8975 33481 9073
rect 33769 8975 33867 9073
rect 34631 8975 34729 9073
rect 35017 8975 35115 9073
rect 35879 8975 35977 9073
rect 36265 8975 36363 9073
rect 37127 8975 37225 9073
rect 37513 8975 37611 9073
rect 38375 8975 38473 9073
rect 38761 8975 38859 9073
rect 39623 8975 39721 9073
rect 40009 8975 40107 9073
rect 40871 8975 40969 9073
rect 41257 8975 41355 9073
rect 42119 8975 42217 9073
rect 42505 8975 42603 9073
rect 43367 8975 43465 9073
rect 43753 8975 43851 9073
rect 44615 8975 44713 9073
rect 45001 8975 45099 9073
rect 45863 8975 45961 9073
rect 46249 8975 46347 9073
rect 47111 8975 47209 9073
rect 47497 8975 47595 9073
rect 48359 8975 48457 9073
rect 48745 8975 48843 9073
rect 49607 8975 49705 9073
rect 49993 8975 50091 9073
rect 50855 8975 50953 9073
rect 51241 8975 51339 9073
rect 52103 8975 52201 9073
rect 52489 8975 52587 9073
rect 53351 8975 53449 9073
rect 11644 8435 11710 8438
rect 11644 8433 32938 8435
rect 11644 8377 11649 8433
rect 11705 8377 32938 8433
rect 11644 8375 32938 8377
rect 11644 8372 11710 8375
rect 13544 8286 13610 8289
rect 0 8284 13610 8286
rect 0 8228 13549 8284
rect 13605 8228 13610 8284
rect 0 8226 13610 8228
rect 13544 8223 13610 8226
rect 6708 7663 6806 7684
rect 6708 7607 6729 7663
rect 6785 7607 6806 7663
rect 6708 7586 6806 7607
rect 14232 7426 14330 7524
rect 15480 7426 15578 7524
rect 16728 7426 16826 7524
rect 17976 7426 18074 7524
rect 19224 7426 19322 7524
rect 20472 7426 20570 7524
rect 21720 7426 21818 7524
rect 22968 7426 23066 7524
rect 24216 7426 24314 7524
rect 25464 7426 25562 7524
rect 26712 7426 26810 7524
rect 27960 7426 28058 7524
rect 29208 7426 29306 7524
rect 30456 7426 30554 7524
rect 31704 7426 31802 7524
rect 32952 7426 33050 7524
rect 34200 7426 34298 7524
rect 35448 7426 35546 7524
rect 36696 7426 36794 7524
rect 37944 7426 38042 7524
rect 39192 7426 39290 7524
rect 40440 7426 40538 7524
rect 41688 7426 41786 7524
rect 42936 7426 43034 7524
rect 44184 7426 44282 7524
rect 45432 7426 45530 7524
rect 46680 7426 46778 7524
rect 47928 7426 48026 7524
rect 49176 7426 49274 7524
rect 50424 7426 50522 7524
rect 51672 7426 51770 7524
rect 52920 7426 53018 7524
rect 7123 6958 7189 6961
rect 7752 6958 7818 6961
rect 7123 6956 7818 6958
rect 7123 6900 7128 6956
rect 7184 6900 7757 6956
rect 7813 6900 7818 6956
rect 7123 6898 7818 6900
rect 7123 6895 7189 6898
rect 7752 6895 7818 6898
rect 7752 6748 7818 6751
rect 7752 6746 12313 6748
rect 7752 6690 7757 6746
rect 7813 6690 12313 6746
rect 7752 6688 12313 6690
rect 7752 6685 7818 6688
rect 7616 6624 7682 6627
rect 7616 6622 12313 6624
rect 7616 6566 7621 6622
rect 7677 6566 12313 6622
rect 7616 6564 12313 6566
rect 7616 6561 7682 6564
rect 6708 6249 6806 6270
rect 6708 6193 6729 6249
rect 6785 6193 6806 6249
rect 6708 6172 6806 6193
rect 11768 5908 11834 5911
rect 11768 5906 32564 5908
rect 11768 5850 11773 5906
rect 11829 5850 32564 5906
rect 11768 5848 32564 5850
rect 11768 5845 11834 5848
rect 14059 5677 14157 5775
rect 15307 5677 15405 5775
rect 16555 5677 16653 5775
rect 17803 5677 17901 5775
rect 19051 5677 19149 5775
rect 20299 5677 20397 5775
rect 21547 5677 21645 5775
rect 22795 5677 22893 5775
rect 24043 5677 24141 5775
rect 25291 5677 25389 5775
rect 26539 5677 26637 5775
rect 27787 5677 27885 5775
rect 29035 5677 29133 5775
rect 30283 5677 30381 5775
rect 31531 5677 31629 5775
rect 32779 5677 32877 5775
rect 34027 5677 34125 5775
rect 35275 5677 35373 5775
rect 36523 5677 36621 5775
rect 37771 5677 37869 5775
rect 39019 5677 39117 5775
rect 40267 5677 40365 5775
rect 41515 5677 41613 5775
rect 42763 5677 42861 5775
rect 44011 5677 44109 5775
rect 45259 5677 45357 5775
rect 46507 5677 46605 5775
rect 47755 5677 47853 5775
rect 49003 5677 49101 5775
rect 50251 5677 50349 5775
rect 51499 5677 51597 5775
rect 52747 5677 52845 5775
rect 7123 5544 7189 5547
rect 7616 5544 7682 5547
rect 7123 5542 7682 5544
rect 7123 5486 7128 5542
rect 7184 5486 7621 5542
rect 7677 5486 7682 5542
rect 7123 5484 7682 5486
rect 7123 5481 7189 5484
rect 7616 5481 7682 5484
rect 13977 4903 14075 5001
rect 15225 4903 15323 5001
rect 16473 4903 16571 5001
rect 17721 4903 17819 5001
rect 18969 4903 19067 5001
rect 20217 4903 20315 5001
rect 21465 4903 21563 5001
rect 22713 4903 22811 5001
rect 23961 4903 24059 5001
rect 25209 4903 25307 5001
rect 26457 4903 26555 5001
rect 27705 4903 27803 5001
rect 28953 4903 29051 5001
rect 30201 4903 30299 5001
rect 31449 4903 31547 5001
rect 32697 4903 32795 5001
rect 33945 4903 34043 5001
rect 35193 4903 35291 5001
rect 36441 4903 36539 5001
rect 37689 4903 37787 5001
rect 38937 4903 39035 5001
rect 40185 4903 40283 5001
rect 41433 4903 41531 5001
rect 42681 4903 42779 5001
rect 43929 4903 44027 5001
rect 45177 4903 45275 5001
rect 46425 4903 46523 5001
rect 47673 4903 47771 5001
rect 48921 4903 49019 5001
rect 50169 4903 50267 5001
rect 51417 4903 51515 5001
rect 52665 4903 52763 5001
rect 6708 4835 6806 4856
rect 6708 4779 6729 4835
rect 6785 4779 6806 4835
rect 6708 4758 6806 4779
rect 13989 4065 14087 4163
rect 15237 4065 15335 4163
rect 16485 4065 16583 4163
rect 17733 4065 17831 4163
rect 18981 4065 19079 4163
rect 20229 4065 20327 4163
rect 21477 4065 21575 4163
rect 22725 4065 22823 4163
rect 23973 4065 24071 4163
rect 25221 4065 25319 4163
rect 26469 4065 26567 4163
rect 27717 4065 27815 4163
rect 28965 4065 29063 4163
rect 30213 4065 30311 4163
rect 31461 4065 31559 4163
rect 32709 4065 32807 4163
rect 33957 4065 34055 4163
rect 35205 4065 35303 4163
rect 36453 4065 36551 4163
rect 37701 4065 37799 4163
rect 38949 4065 39047 4163
rect 40197 4065 40295 4163
rect 41445 4065 41543 4163
rect 42693 4065 42791 4163
rect 43941 4065 44039 4163
rect 45189 4065 45287 4163
rect 46437 4065 46535 4163
rect 47685 4065 47783 4163
rect 48933 4065 49031 4163
rect 50181 4065 50279 4163
rect 51429 4065 51527 4163
rect 52677 4065 52775 4163
rect 13989 3743 14087 3841
rect 15237 3743 15335 3841
rect 16485 3743 16583 3841
rect 17733 3743 17831 3841
rect 18981 3743 19079 3841
rect 20229 3743 20327 3841
rect 21477 3743 21575 3841
rect 22725 3743 22823 3841
rect 23973 3743 24071 3841
rect 25221 3743 25319 3841
rect 26469 3743 26567 3841
rect 27717 3743 27815 3841
rect 28965 3743 29063 3841
rect 30213 3743 30311 3841
rect 31461 3743 31559 3841
rect 32709 3743 32807 3841
rect 33957 3743 34055 3841
rect 35205 3743 35303 3841
rect 36453 3743 36551 3841
rect 37701 3743 37799 3841
rect 38949 3743 39047 3841
rect 40197 3743 40295 3841
rect 41445 3743 41543 3841
rect 42693 3743 42791 3841
rect 43941 3743 44039 3841
rect 45189 3743 45287 3841
rect 46437 3743 46535 3841
rect 47685 3743 47783 3841
rect 48933 3743 49031 3841
rect 50181 3743 50279 3841
rect 51429 3743 51527 3841
rect 52677 3743 52775 3841
rect 13875 2950 13973 3048
rect 15123 2950 15221 3048
rect 16371 2950 16469 3048
rect 17619 2950 17717 3048
rect 18867 2950 18965 3048
rect 20115 2950 20213 3048
rect 21363 2950 21461 3048
rect 22611 2950 22709 3048
rect 23859 2950 23957 3048
rect 25107 2950 25205 3048
rect 26355 2950 26453 3048
rect 27603 2950 27701 3048
rect 28851 2950 28949 3048
rect 30099 2950 30197 3048
rect 31347 2950 31445 3048
rect 32595 2950 32693 3048
rect 33843 2950 33941 3048
rect 35091 2950 35189 3048
rect 36339 2950 36437 3048
rect 37587 2950 37685 3048
rect 38835 2950 38933 3048
rect 40083 2950 40181 3048
rect 41331 2950 41429 3048
rect 42579 2950 42677 3048
rect 43827 2950 43925 3048
rect 45075 2950 45173 3048
rect 46323 2950 46421 3048
rect 47571 2950 47669 3048
rect 48819 2950 48917 3048
rect 50067 2950 50165 3048
rect 51315 2950 51413 3048
rect 52563 2950 52661 3048
rect 13864 2513 13962 2611
rect 15112 2513 15210 2611
rect 16360 2513 16458 2611
rect 17608 2513 17706 2611
rect 18856 2513 18954 2611
rect 20104 2513 20202 2611
rect 21352 2513 21450 2611
rect 22600 2513 22698 2611
rect 23848 2513 23946 2611
rect 25096 2513 25194 2611
rect 26344 2513 26442 2611
rect 27592 2513 27690 2611
rect 28840 2513 28938 2611
rect 30088 2513 30186 2611
rect 31336 2513 31434 2611
rect 32584 2513 32682 2611
rect 33832 2513 33930 2611
rect 35080 2513 35178 2611
rect 36328 2513 36426 2611
rect 37576 2513 37674 2611
rect 38824 2513 38922 2611
rect 40072 2513 40170 2611
rect 41320 2513 41418 2611
rect 42568 2513 42666 2611
rect 43816 2513 43914 2611
rect 45064 2513 45162 2611
rect 46312 2513 46410 2611
rect 47560 2513 47658 2611
rect 48808 2513 48906 2611
rect 50056 2513 50154 2611
rect 51304 2513 51402 2611
rect 52552 2513 52650 2611
rect 13985 2181 14083 2279
rect 15233 2181 15331 2279
rect 16481 2181 16579 2279
rect 17729 2181 17827 2279
rect 18977 2181 19075 2279
rect 20225 2181 20323 2279
rect 21473 2181 21571 2279
rect 22721 2181 22819 2279
rect 23969 2181 24067 2279
rect 25217 2181 25315 2279
rect 26465 2181 26563 2279
rect 27713 2181 27811 2279
rect 28961 2181 29059 2279
rect 30209 2181 30307 2279
rect 31457 2181 31555 2279
rect 32705 2181 32803 2279
rect 33953 2181 34051 2279
rect 35201 2181 35299 2279
rect 36449 2181 36547 2279
rect 37697 2181 37795 2279
rect 38945 2181 39043 2279
rect 40193 2181 40291 2279
rect 41441 2181 41539 2279
rect 42689 2181 42787 2279
rect 43937 2181 44035 2279
rect 45185 2181 45283 2279
rect 46433 2181 46531 2279
rect 47681 2181 47779 2279
rect 48929 2181 49027 2279
rect 50177 2181 50275 2279
rect 51425 2181 51523 2279
rect 52673 2181 52771 2279
rect 13870 1979 13968 2077
rect 15118 1979 15216 2077
rect 16366 1979 16464 2077
rect 17614 1979 17712 2077
rect 18862 1979 18960 2077
rect 20110 1979 20208 2077
rect 21358 1979 21456 2077
rect 22606 1979 22704 2077
rect 23854 1979 23952 2077
rect 25102 1979 25200 2077
rect 26350 1979 26448 2077
rect 27598 1979 27696 2077
rect 28846 1979 28944 2077
rect 30094 1979 30192 2077
rect 31342 1979 31440 2077
rect 32590 1979 32688 2077
rect 33838 1979 33936 2077
rect 35086 1979 35184 2077
rect 36334 1979 36432 2077
rect 37582 1979 37680 2077
rect 38830 1979 38928 2077
rect 40078 1979 40176 2077
rect 41326 1979 41424 2077
rect 42574 1979 42672 2077
rect 43822 1979 43920 2077
rect 45070 1979 45168 2077
rect 46318 1979 46416 2077
rect 47566 1979 47664 2077
rect 48814 1979 48912 2077
rect 50062 1979 50160 2077
rect 51310 1979 51408 2077
rect 52558 1979 52656 2077
rect 13884 1563 13982 1661
rect 15132 1563 15230 1661
rect 16380 1563 16478 1661
rect 17628 1563 17726 1661
rect 18876 1563 18974 1661
rect 20124 1563 20222 1661
rect 21372 1563 21470 1661
rect 22620 1563 22718 1661
rect 23868 1563 23966 1661
rect 25116 1563 25214 1661
rect 26364 1563 26462 1661
rect 27612 1563 27710 1661
rect 28860 1563 28958 1661
rect 30108 1563 30206 1661
rect 31356 1563 31454 1661
rect 32604 1563 32702 1661
rect 33852 1563 33950 1661
rect 35100 1563 35198 1661
rect 36348 1563 36446 1661
rect 37596 1563 37694 1661
rect 38844 1563 38942 1661
rect 40092 1563 40190 1661
rect 41340 1563 41438 1661
rect 42588 1563 42686 1661
rect 43836 1563 43934 1661
rect 45084 1563 45182 1661
rect 46332 1563 46430 1661
rect 47580 1563 47678 1661
rect 48828 1563 48926 1661
rect 50076 1563 50174 1661
rect 51324 1563 51422 1661
rect 52572 1563 52670 1661
rect 12234 1120 12332 1218
rect 53544 1120 53642 1218
rect 11892 597 11958 600
rect 11892 595 32938 597
rect 11892 539 11897 595
rect 11953 539 32938 595
rect 11892 537 32938 539
rect 11892 534 11958 537
rect 12234 0 12332 98
rect 53544 0 53642 98
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_0
timestamp 1636140361
transform 1 0 55062 0 1 13424
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_0
timestamp 1636140361
transform 1 0 55065 0 1 13423
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_1
timestamp 1636140361
transform 1 0 55062 0 1 13184
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_1
timestamp 1636140361
transform 1 0 55065 0 1 13183
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_2
timestamp 1636140361
transform 1 0 55062 0 1 12634
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_2
timestamp 1636140361
transform 1 0 55065 0 1 12633
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_3
timestamp 1636140361
transform 1 0 55062 0 1 12394
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_3
timestamp 1636140361
transform 1 0 55065 0 1 12393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_4
timestamp 1636140361
transform 1 0 55062 0 1 11844
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_4
timestamp 1636140361
transform 1 0 55065 0 1 11843
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_5
timestamp 1636140361
transform 1 0 55062 0 1 11604
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_5
timestamp 1636140361
transform 1 0 55065 0 1 11603
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_6
timestamp 1636140361
transform 1 0 55062 0 1 11054
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_6
timestamp 1636140361
transform 1 0 55065 0 1 11053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_7
timestamp 1636140361
transform 1 0 55062 0 1 10814
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_7
timestamp 1636140361
transform 1 0 55065 0 1 10813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_8
timestamp 1636140361
transform 1 0 55062 0 1 10264
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_8
timestamp 1636140361
transform 1 0 55065 0 1 10263
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_9
timestamp 1636140361
transform 1 0 55062 0 1 16584
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_9
timestamp 1636140361
transform 1 0 55065 0 1 16583
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_10
timestamp 1636140361
transform 1 0 55062 0 1 16344
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_10
timestamp 1636140361
transform 1 0 55065 0 1 16343
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_11
timestamp 1636140361
transform 1 0 55062 0 1 15794
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_11
timestamp 1636140361
transform 1 0 55065 0 1 15793
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_12
timestamp 1636140361
transform 1 0 55062 0 1 15554
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_12
timestamp 1636140361
transform 1 0 55065 0 1 15553
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_13
timestamp 1636140361
transform 1 0 55062 0 1 15004
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_13
timestamp 1636140361
transform 1 0 55065 0 1 15003
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_14
timestamp 1636140361
transform 1 0 55062 0 1 14764
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_14
timestamp 1636140361
transform 1 0 55065 0 1 14763
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_15
timestamp 1636140361
transform 1 0 55062 0 1 14214
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_15
timestamp 1636140361
transform 1 0 55065 0 1 14213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_16
timestamp 1636140361
transform 1 0 55062 0 1 13974
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_16
timestamp 1636140361
transform 1 0 55065 0 1 13973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_17
timestamp 1636140361
transform 1 0 55062 0 1 20294
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_17
timestamp 1636140361
transform 1 0 55065 0 1 20293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_18
timestamp 1636140361
transform 1 0 55062 0 1 19744
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_18
timestamp 1636140361
transform 1 0 55065 0 1 19743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_19
timestamp 1636140361
transform 1 0 55062 0 1 19504
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_19
timestamp 1636140361
transform 1 0 55065 0 1 19503
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_20
timestamp 1636140361
transform 1 0 55062 0 1 18954
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_20
timestamp 1636140361
transform 1 0 55065 0 1 18953
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_21
timestamp 1636140361
transform 1 0 55062 0 1 18714
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_21
timestamp 1636140361
transform 1 0 55065 0 1 18713
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_22
timestamp 1636140361
transform 1 0 55062 0 1 18164
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_22
timestamp 1636140361
transform 1 0 55065 0 1 18163
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_23
timestamp 1636140361
transform 1 0 55062 0 1 17924
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_23
timestamp 1636140361
transform 1 0 55065 0 1 17923
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_24
timestamp 1636140361
transform 1 0 55062 0 1 17374
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_24
timestamp 1636140361
transform 1 0 55065 0 1 17373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_25
timestamp 1636140361
transform 1 0 55062 0 1 17134
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_25
timestamp 1636140361
transform 1 0 55065 0 1 17133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_26
timestamp 1636140361
transform 1 0 55062 0 1 33174
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_26
timestamp 1636140361
transform 1 0 55065 0 1 33173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_27
timestamp 1636140361
transform 1 0 55062 0 1 32934
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_27
timestamp 1636140361
transform 1 0 55065 0 1 32933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_28
timestamp 1636140361
transform 1 0 55062 0 1 32384
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_28
timestamp 1636140361
transform 1 0 55065 0 1 32383
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_29
timestamp 1636140361
transform 1 0 55062 0 1 32144
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_29
timestamp 1636140361
transform 1 0 55065 0 1 32143
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_30
timestamp 1636140361
transform 1 0 55062 0 1 31594
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_30
timestamp 1636140361
transform 1 0 55065 0 1 31593
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_31
timestamp 1636140361
transform 1 0 55062 0 1 31354
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_31
timestamp 1636140361
transform 1 0 55065 0 1 31353
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_32
timestamp 1636140361
transform 1 0 55062 0 1 30804
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_32
timestamp 1636140361
transform 1 0 55065 0 1 30803
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_33
timestamp 1636140361
transform 1 0 55062 0 1 30564
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_33
timestamp 1636140361
transform 1 0 55065 0 1 30563
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_34
timestamp 1636140361
transform 1 0 55062 0 1 30014
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_34
timestamp 1636140361
transform 1 0 55065 0 1 30013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_35
timestamp 1636140361
transform 1 0 55062 0 1 29774
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_35
timestamp 1636140361
transform 1 0 55065 0 1 29773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_36
timestamp 1636140361
transform 1 0 55062 0 1 29224
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_36
timestamp 1636140361
transform 1 0 55065 0 1 29223
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_37
timestamp 1636140361
transform 1 0 55062 0 1 28984
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_37
timestamp 1636140361
transform 1 0 55065 0 1 28983
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_38
timestamp 1636140361
transform 1 0 55062 0 1 28434
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_38
timestamp 1636140361
transform 1 0 55065 0 1 28433
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_39
timestamp 1636140361
transform 1 0 55062 0 1 28194
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_39
timestamp 1636140361
transform 1 0 55065 0 1 28193
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_40
timestamp 1636140361
transform 1 0 55062 0 1 27644
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_40
timestamp 1636140361
transform 1 0 55065 0 1 27643
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_41
timestamp 1636140361
transform 1 0 55062 0 1 27404
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_41
timestamp 1636140361
transform 1 0 55065 0 1 27403
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_42
timestamp 1636140361
transform 1 0 55062 0 1 26854
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_42
timestamp 1636140361
transform 1 0 55065 0 1 26853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_43
timestamp 1636140361
transform 1 0 55062 0 1 26614
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_43
timestamp 1636140361
transform 1 0 55065 0 1 26613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_44
timestamp 1636140361
transform 1 0 55062 0 1 26064
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_44
timestamp 1636140361
transform 1 0 55065 0 1 26063
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_45
timestamp 1636140361
transform 1 0 55062 0 1 25824
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_45
timestamp 1636140361
transform 1 0 55065 0 1 25823
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_46
timestamp 1636140361
transform 1 0 55062 0 1 25274
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_46
timestamp 1636140361
transform 1 0 55065 0 1 25273
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_47
timestamp 1636140361
transform 1 0 55062 0 1 25034
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_47
timestamp 1636140361
transform 1 0 55065 0 1 25033
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_48
timestamp 1636140361
transform 1 0 55062 0 1 24484
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_48
timestamp 1636140361
transform 1 0 55065 0 1 24483
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_49
timestamp 1636140361
transform 1 0 55062 0 1 24244
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_49
timestamp 1636140361
transform 1 0 55065 0 1 24243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_50
timestamp 1636140361
transform 1 0 55062 0 1 23694
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_50
timestamp 1636140361
transform 1 0 55065 0 1 23693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_51
timestamp 1636140361
transform 1 0 55062 0 1 23454
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_51
timestamp 1636140361
transform 1 0 55065 0 1 23453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_52
timestamp 1636140361
transform 1 0 55062 0 1 22904
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_52
timestamp 1636140361
transform 1 0 55065 0 1 22903
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_53
timestamp 1636140361
transform 1 0 55062 0 1 22664
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_53
timestamp 1636140361
transform 1 0 55065 0 1 22663
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_54
timestamp 1636140361
transform 1 0 55062 0 1 22114
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_54
timestamp 1636140361
transform 1 0 55065 0 1 22113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_55
timestamp 1636140361
transform 1 0 55062 0 1 21874
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_55
timestamp 1636140361
transform 1 0 55065 0 1 21873
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_56
timestamp 1636140361
transform 1 0 55062 0 1 21324
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_56
timestamp 1636140361
transform 1 0 55065 0 1 21323
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_57
timestamp 1636140361
transform 1 0 55062 0 1 21084
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_57
timestamp 1636140361
transform 1 0 55065 0 1 21083
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_58
timestamp 1636140361
transform 1 0 55062 0 1 20534
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_58
timestamp 1636140361
transform 1 0 55065 0 1 20533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_59
timestamp 1636140361
transform 1 0 12124 0 1 10814
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_59
timestamp 1636140361
transform 1 0 12127 0 1 10813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_60
timestamp 1636140361
transform 1 0 12124 0 1 10264
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_60
timestamp 1636140361
transform 1 0 12127 0 1 10263
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_0
timestamp 1636140361
transform 1 0 13544 0 1 8219
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_61
timestamp 1636140361
transform 1 0 13545 0 1 8224
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf  sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf_0
timestamp 1636140361
transform 1 0 5989 0 1 4790
box -36 0 1536 2862
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_62
timestamp 1636140361
transform 1 0 12124 0 1 16584
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_61
timestamp 1636140361
transform 1 0 12127 0 1 16583
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_1
timestamp 1636140361
transform 1 0 6724 0 1 7598
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_63
timestamp 1636140361
transform 1 0 6725 0 1 7603
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_62
timestamp 1636140361
transform 1 0 6728 0 1 7602
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_2
timestamp 1636140361
transform 1 0 6724 0 1 4770
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_64
timestamp 1636140361
transform 1 0 6725 0 1 4775
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_63
timestamp 1636140361
transform 1 0 6728 0 1 4774
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_3
timestamp 1636140361
transform 1 0 6724 0 1 6184
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_65
timestamp 1636140361
transform 1 0 6725 0 1 6189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_64
timestamp 1636140361
transform 1 0 6728 0 1 6188
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_66
timestamp 1636140361
transform 1 0 12124 0 1 16344
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_65
timestamp 1636140361
transform 1 0 12127 0 1 16343
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_67
timestamp 1636140361
transform 1 0 12124 0 1 15794
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_66
timestamp 1636140361
transform 1 0 12127 0 1 15793
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_68
timestamp 1636140361
transform 1 0 12124 0 1 15554
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_67
timestamp 1636140361
transform 1 0 12127 0 1 15553
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_69
timestamp 1636140361
transform 1 0 12124 0 1 15004
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_68
timestamp 1636140361
transform 1 0 12127 0 1 15003
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_70
timestamp 1636140361
transform 1 0 12124 0 1 14764
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_69
timestamp 1636140361
transform 1 0 12127 0 1 14763
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_71
timestamp 1636140361
transform 1 0 12124 0 1 14214
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_70
timestamp 1636140361
transform 1 0 12127 0 1 14213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_72
timestamp 1636140361
transform 1 0 12124 0 1 13974
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_71
timestamp 1636140361
transform 1 0 12127 0 1 13973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_73
timestamp 1636140361
transform 1 0 12124 0 1 13424
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_72
timestamp 1636140361
transform 1 0 12127 0 1 13423
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_74
timestamp 1636140361
transform 1 0 12124 0 1 13184
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_73
timestamp 1636140361
transform 1 0 12127 0 1 13183
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_4
timestamp 1636140361
transform 1 0 11768 0 1 5841
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_5
timestamp 1636140361
transform 1 0 11892 0 1 530
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_6
timestamp 1636140361
transform 1 0 11644 0 1 8368
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_7
timestamp 1636140361
transform 1 0 7752 0 1 6681
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_8
timestamp 1636140361
transform 1 0 7123 0 1 6891
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_75
timestamp 1636140361
transform 1 0 7124 0 1 6896
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_74
timestamp 1636140361
transform 1 0 7127 0 1 6895
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_9
timestamp 1636140361
transform 1 0 7752 0 1 6891
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_10
timestamp 1636140361
transform 1 0 7616 0 1 6557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_11
timestamp 1636140361
transform 1 0 7123 0 1 5477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_76
timestamp 1636140361
transform 1 0 7124 0 1 5482
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_75
timestamp 1636140361
transform 1 0 7127 0 1 5481
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_12
timestamp 1636140361
transform 1 0 7616 0 1 5477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_77
timestamp 1636140361
transform 1 0 12124 0 1 10024
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_76
timestamp 1636140361
transform 1 0 12127 0 1 10023
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_78
timestamp 1636140361
transform 1 0 12124 0 1 12634
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_77
timestamp 1636140361
transform 1 0 12127 0 1 12633
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_79
timestamp 1636140361
transform 1 0 12124 0 1 12394
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_78
timestamp 1636140361
transform 1 0 12127 0 1 12393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_80
timestamp 1636140361
transform 1 0 12124 0 1 11844
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_79
timestamp 1636140361
transform 1 0 12127 0 1 11843
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_81
timestamp 1636140361
transform 1 0 12124 0 1 11604
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_80
timestamp 1636140361
transform 1 0 12127 0 1 11603
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_82
timestamp 1636140361
transform 1 0 12124 0 1 11054
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_81
timestamp 1636140361
transform 1 0 12127 0 1 11053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_82
timestamp 1636140361
transform 1 0 12127 0 1 18163
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_83
timestamp 1636140361
transform 1 0 12124 0 1 17924
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_83
timestamp 1636140361
transform 1 0 12127 0 1 17923
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_84
timestamp 1636140361
transform 1 0 12124 0 1 17374
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_84
timestamp 1636140361
transform 1 0 12127 0 1 17373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_85
timestamp 1636140361
transform 1 0 12124 0 1 17134
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_85
timestamp 1636140361
transform 1 0 12127 0 1 17133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_86
timestamp 1636140361
transform 1 0 12124 0 1 33174
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_86
timestamp 1636140361
transform 1 0 12127 0 1 33173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_87
timestamp 1636140361
transform 1 0 12124 0 1 32934
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_87
timestamp 1636140361
transform 1 0 12127 0 1 32933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_88
timestamp 1636140361
transform 1 0 12124 0 1 32384
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_88
timestamp 1636140361
transform 1 0 12127 0 1 32383
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_89
timestamp 1636140361
transform 1 0 12124 0 1 32144
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_89
timestamp 1636140361
transform 1 0 12127 0 1 32143
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_90
timestamp 1636140361
transform 1 0 12124 0 1 31594
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_90
timestamp 1636140361
transform 1 0 12127 0 1 31593
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_91
timestamp 1636140361
transform 1 0 12124 0 1 31354
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_91
timestamp 1636140361
transform 1 0 12127 0 1 31353
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_92
timestamp 1636140361
transform 1 0 12124 0 1 30804
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_92
timestamp 1636140361
transform 1 0 12127 0 1 30803
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_93
timestamp 1636140361
transform 1 0 12124 0 1 30564
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_93
timestamp 1636140361
transform 1 0 12127 0 1 30563
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_94
timestamp 1636140361
transform 1 0 12124 0 1 30014
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_94
timestamp 1636140361
transform 1 0 12127 0 1 30013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_95
timestamp 1636140361
transform 1 0 12124 0 1 29774
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_95
timestamp 1636140361
transform 1 0 12127 0 1 29773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_96
timestamp 1636140361
transform 1 0 12124 0 1 29224
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_96
timestamp 1636140361
transform 1 0 12127 0 1 29223
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_97
timestamp 1636140361
transform 1 0 12124 0 1 28984
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_97
timestamp 1636140361
transform 1 0 12127 0 1 28983
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_98
timestamp 1636140361
transform 1 0 12124 0 1 28434
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_98
timestamp 1636140361
transform 1 0 12127 0 1 28433
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_99
timestamp 1636140361
transform 1 0 12124 0 1 28194
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_99
timestamp 1636140361
transform 1 0 12127 0 1 28193
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_100
timestamp 1636140361
transform 1 0 12124 0 1 27644
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_100
timestamp 1636140361
transform 1 0 12127 0 1 27643
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_101
timestamp 1636140361
transform 1 0 12124 0 1 27404
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_101
timestamp 1636140361
transform 1 0 12127 0 1 27403
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_102
timestamp 1636140361
transform 1 0 12124 0 1 26854
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_102
timestamp 1636140361
transform 1 0 12127 0 1 26853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_103
timestamp 1636140361
transform 1 0 12124 0 1 26614
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_103
timestamp 1636140361
transform 1 0 12127 0 1 26613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_104
timestamp 1636140361
transform 1 0 12124 0 1 26064
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_104
timestamp 1636140361
transform 1 0 12127 0 1 26063
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_105
timestamp 1636140361
transform 1 0 12124 0 1 25824
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_105
timestamp 1636140361
transform 1 0 12127 0 1 25823
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_106
timestamp 1636140361
transform 1 0 12124 0 1 25274
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_106
timestamp 1636140361
transform 1 0 12127 0 1 25273
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_107
timestamp 1636140361
transform 1 0 12124 0 1 25034
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_107
timestamp 1636140361
transform 1 0 12127 0 1 25033
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_108
timestamp 1636140361
transform 1 0 12124 0 1 24484
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_108
timestamp 1636140361
transform 1 0 12127 0 1 24483
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_109
timestamp 1636140361
transform 1 0 12124 0 1 24244
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_109
timestamp 1636140361
transform 1 0 12127 0 1 24243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_110
timestamp 1636140361
transform 1 0 12124 0 1 23694
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_110
timestamp 1636140361
transform 1 0 12127 0 1 23693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_111
timestamp 1636140361
transform 1 0 12124 0 1 23454
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_111
timestamp 1636140361
transform 1 0 12127 0 1 23453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_112
timestamp 1636140361
transform 1 0 12124 0 1 22904
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_112
timestamp 1636140361
transform 1 0 12127 0 1 22903
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_113
timestamp 1636140361
transform 1 0 12124 0 1 22664
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_113
timestamp 1636140361
transform 1 0 12127 0 1 22663
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_114
timestamp 1636140361
transform 1 0 12124 0 1 22114
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_114
timestamp 1636140361
transform 1 0 12127 0 1 22113
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_115
timestamp 1636140361
transform 1 0 12124 0 1 21874
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_115
timestamp 1636140361
transform 1 0 12127 0 1 21873
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_116
timestamp 1636140361
transform 1 0 12124 0 1 21324
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_116
timestamp 1636140361
transform 1 0 12127 0 1 21323
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_117
timestamp 1636140361
transform 1 0 12124 0 1 21084
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_117
timestamp 1636140361
transform 1 0 12127 0 1 21083
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_118
timestamp 1636140361
transform 1 0 12124 0 1 20534
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_118
timestamp 1636140361
transform 1 0 12127 0 1 20533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_119
timestamp 1636140361
transform 1 0 12124 0 1 20294
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_119
timestamp 1636140361
transform 1 0 12127 0 1 20293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_120
timestamp 1636140361
transform 1 0 12124 0 1 19744
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_120
timestamp 1636140361
transform 1 0 12127 0 1 19743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_121
timestamp 1636140361
transform 1 0 12124 0 1 19504
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_121
timestamp 1636140361
transform 1 0 12127 0 1 19503
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_122
timestamp 1636140361
transform 1 0 12124 0 1 18954
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_122
timestamp 1636140361
transform 1 0 12127 0 1 18953
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_123
timestamp 1636140361
transform 1 0 12124 0 1 18714
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_123
timestamp 1636140361
transform 1 0 12127 0 1 18713
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_124
timestamp 1636140361
transform 1 0 12124 0 1 18164
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_124
timestamp 1636140361
transform 1 0 12127 0 1 38463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_125
timestamp 1636140361
transform 1 0 12124 0 1 37914
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_125
timestamp 1636140361
transform 1 0 12127 0 1 37913
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_126
timestamp 1636140361
transform 1 0 12124 0 1 37674
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_126
timestamp 1636140361
transform 1 0 12127 0 1 37673
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_127
timestamp 1636140361
transform 1 0 12124 0 1 37124
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_127
timestamp 1636140361
transform 1 0 12127 0 1 37123
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_128
timestamp 1636140361
transform 1 0 12124 0 1 36884
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_128
timestamp 1636140361
transform 1 0 12127 0 1 36883
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_129
timestamp 1636140361
transform 1 0 12124 0 1 36334
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_129
timestamp 1636140361
transform 1 0 12127 0 1 36333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_130
timestamp 1636140361
transform 1 0 12124 0 1 36094
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_130
timestamp 1636140361
transform 1 0 12127 0 1 36093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_131
timestamp 1636140361
transform 1 0 12124 0 1 35544
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_131
timestamp 1636140361
transform 1 0 12127 0 1 35543
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_132
timestamp 1636140361
transform 1 0 12124 0 1 35304
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_132
timestamp 1636140361
transform 1 0 12127 0 1 35303
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_133
timestamp 1636140361
transform 1 0 12124 0 1 34754
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_133
timestamp 1636140361
transform 1 0 12127 0 1 34753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_134
timestamp 1636140361
transform 1 0 12124 0 1 34514
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_134
timestamp 1636140361
transform 1 0 12127 0 1 34513
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_135
timestamp 1636140361
transform 1 0 12124 0 1 33964
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_135
timestamp 1636140361
transform 1 0 12127 0 1 33963
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_136
timestamp 1636140361
transform 1 0 12124 0 1 33724
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_136
timestamp 1636140361
transform 1 0 12127 0 1 33723
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_137
timestamp 1636140361
transform 1 0 12127 0 1 48733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_137
timestamp 1636140361
transform 1 0 12124 0 1 48184
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_138
timestamp 1636140361
transform 1 0 12127 0 1 48183
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_138
timestamp 1636140361
transform 1 0 12124 0 1 47944
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_139
timestamp 1636140361
transform 1 0 12127 0 1 47943
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_139
timestamp 1636140361
transform 1 0 12124 0 1 47394
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_140
timestamp 1636140361
transform 1 0 12127 0 1 47393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_140
timestamp 1636140361
transform 1 0 12124 0 1 47154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_141
timestamp 1636140361
transform 1 0 12127 0 1 47153
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_141
timestamp 1636140361
transform 1 0 12124 0 1 46604
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_142
timestamp 1636140361
transform 1 0 12127 0 1 46603
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_142
timestamp 1636140361
transform 1 0 12124 0 1 46364
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_143
timestamp 1636140361
transform 1 0 12127 0 1 46363
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_143
timestamp 1636140361
transform 1 0 12124 0 1 45814
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_144
timestamp 1636140361
transform 1 0 12127 0 1 45813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_144
timestamp 1636140361
transform 1 0 12124 0 1 45574
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_145
timestamp 1636140361
transform 1 0 12127 0 1 45573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_145
timestamp 1636140361
transform 1 0 12124 0 1 45024
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_146
timestamp 1636140361
transform 1 0 12127 0 1 45023
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_146
timestamp 1636140361
transform 1 0 12124 0 1 44784
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_147
timestamp 1636140361
transform 1 0 12127 0 1 44783
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_147
timestamp 1636140361
transform 1 0 12124 0 1 44234
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_148
timestamp 1636140361
transform 1 0 12127 0 1 44233
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_148
timestamp 1636140361
transform 1 0 12124 0 1 43994
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_149
timestamp 1636140361
transform 1 0 12127 0 1 43993
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_149
timestamp 1636140361
transform 1 0 12124 0 1 43444
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_150
timestamp 1636140361
transform 1 0 12127 0 1 43443
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_150
timestamp 1636140361
transform 1 0 12124 0 1 43204
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_151
timestamp 1636140361
transform 1 0 12127 0 1 43203
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_151
timestamp 1636140361
transform 1 0 12124 0 1 42654
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_152
timestamp 1636140361
transform 1 0 12127 0 1 42653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_152
timestamp 1636140361
transform 1 0 12124 0 1 42414
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_153
timestamp 1636140361
transform 1 0 12127 0 1 42413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_153
timestamp 1636140361
transform 1 0 12124 0 1 41864
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_154
timestamp 1636140361
transform 1 0 12127 0 1 41863
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_154
timestamp 1636140361
transform 1 0 12124 0 1 41624
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_155
timestamp 1636140361
transform 1 0 12127 0 1 41623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_155
timestamp 1636140361
transform 1 0 12124 0 1 41074
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_156
timestamp 1636140361
transform 1 0 12127 0 1 41073
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_156
timestamp 1636140361
transform 1 0 12124 0 1 40834
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_157
timestamp 1636140361
transform 1 0 12127 0 1 40833
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_157
timestamp 1636140361
transform 1 0 12124 0 1 40284
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_158
timestamp 1636140361
transform 1 0 12127 0 1 40283
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_158
timestamp 1636140361
transform 1 0 12124 0 1 40044
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_159
timestamp 1636140361
transform 1 0 12127 0 1 40043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_159
timestamp 1636140361
transform 1 0 12124 0 1 39494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_160
timestamp 1636140361
transform 1 0 12127 0 1 39493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_160
timestamp 1636140361
transform 1 0 12124 0 1 39254
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_161
timestamp 1636140361
transform 1 0 12127 0 1 39253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_161
timestamp 1636140361
transform 1 0 12124 0 1 38704
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_162
timestamp 1636140361
transform 1 0 12127 0 1 38703
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_162
timestamp 1636140361
transform 1 0 12124 0 1 38464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_163
timestamp 1636140361
transform 1 0 12124 0 1 50314
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_163
timestamp 1636140361
transform 1 0 12127 0 1 50313
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_164
timestamp 1636140361
transform 1 0 12124 0 1 49764
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_164
timestamp 1636140361
transform 1 0 12127 0 1 49763
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_165
timestamp 1636140361
transform 1 0 12124 0 1 49524
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_165
timestamp 1636140361
transform 1 0 12127 0 1 49523
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_166
timestamp 1636140361
transform 1 0 12124 0 1 48974
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_166
timestamp 1636140361
transform 1 0 12127 0 1 48973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_167
timestamp 1636140361
transform 1 0 12124 0 1 48734
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_168
timestamp 1636140361
transform 1 0 12124 0 1 60584
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_167
timestamp 1636140361
transform 1 0 12127 0 1 60583
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_169
timestamp 1636140361
transform 1 0 12124 0 1 60034
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_168
timestamp 1636140361
transform 1 0 12127 0 1 60033
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_170
timestamp 1636140361
transform 1 0 12124 0 1 59794
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_169
timestamp 1636140361
transform 1 0 12127 0 1 59793
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_171
timestamp 1636140361
transform 1 0 12124 0 1 59244
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_170
timestamp 1636140361
transform 1 0 12127 0 1 59243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_172
timestamp 1636140361
transform 1 0 12124 0 1 59004
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_171
timestamp 1636140361
transform 1 0 12127 0 1 59003
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_173
timestamp 1636140361
transform 1 0 12124 0 1 58454
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_172
timestamp 1636140361
transform 1 0 12127 0 1 58453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_174
timestamp 1636140361
transform 1 0 12124 0 1 58214
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_173
timestamp 1636140361
transform 1 0 12127 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_175
timestamp 1636140361
transform 1 0 12124 0 1 57664
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_174
timestamp 1636140361
transform 1 0 12127 0 1 57663
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_176
timestamp 1636140361
transform 1 0 12124 0 1 57424
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_175
timestamp 1636140361
transform 1 0 12127 0 1 57423
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_177
timestamp 1636140361
transform 1 0 12124 0 1 56874
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_176
timestamp 1636140361
transform 1 0 12127 0 1 56873
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_178
timestamp 1636140361
transform 1 0 12124 0 1 56634
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_177
timestamp 1636140361
transform 1 0 12127 0 1 56633
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_179
timestamp 1636140361
transform 1 0 12124 0 1 56084
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_178
timestamp 1636140361
transform 1 0 12127 0 1 56083
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_180
timestamp 1636140361
transform 1 0 12124 0 1 55844
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_179
timestamp 1636140361
transform 1 0 12127 0 1 55843
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_181
timestamp 1636140361
transform 1 0 12124 0 1 55294
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_180
timestamp 1636140361
transform 1 0 12127 0 1 55293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_182
timestamp 1636140361
transform 1 0 12124 0 1 55054
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_181
timestamp 1636140361
transform 1 0 12127 0 1 55053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_183
timestamp 1636140361
transform 1 0 12124 0 1 54504
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_182
timestamp 1636140361
transform 1 0 12127 0 1 54503
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_184
timestamp 1636140361
transform 1 0 12124 0 1 54264
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_183
timestamp 1636140361
transform 1 0 12127 0 1 54263
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_185
timestamp 1636140361
transform 1 0 12124 0 1 53714
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_184
timestamp 1636140361
transform 1 0 12127 0 1 53713
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_186
timestamp 1636140361
transform 1 0 12124 0 1 53474
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_185
timestamp 1636140361
transform 1 0 12127 0 1 53473
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_187
timestamp 1636140361
transform 1 0 12124 0 1 52924
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_186
timestamp 1636140361
transform 1 0 12127 0 1 52923
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_188
timestamp 1636140361
transform 1 0 12124 0 1 52684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_187
timestamp 1636140361
transform 1 0 12127 0 1 52683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_189
timestamp 1636140361
transform 1 0 12124 0 1 52134
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_188
timestamp 1636140361
transform 1 0 12127 0 1 52133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_190
timestamp 1636140361
transform 1 0 12124 0 1 51894
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_189
timestamp 1636140361
transform 1 0 12127 0 1 51893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_191
timestamp 1636140361
transform 1 0 12124 0 1 51344
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_190
timestamp 1636140361
transform 1 0 12127 0 1 51343
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_192
timestamp 1636140361
transform 1 0 12124 0 1 51104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_191
timestamp 1636140361
transform 1 0 12127 0 1 51103
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_193
timestamp 1636140361
transform 1 0 12124 0 1 50554
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_192
timestamp 1636140361
transform 1 0 12127 0 1 50553
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_193
timestamp 1636140361
transform 1 0 55065 0 1 48183
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_194
timestamp 1636140361
transform 1 0 55062 0 1 47944
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_194
timestamp 1636140361
transform 1 0 55065 0 1 47943
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_195
timestamp 1636140361
transform 1 0 55062 0 1 47394
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_195
timestamp 1636140361
transform 1 0 55065 0 1 47393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_196
timestamp 1636140361
transform 1 0 55062 0 1 47154
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_196
timestamp 1636140361
transform 1 0 55065 0 1 47153
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_197
timestamp 1636140361
transform 1 0 55062 0 1 46604
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_197
timestamp 1636140361
transform 1 0 55065 0 1 46603
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_198
timestamp 1636140361
transform 1 0 55062 0 1 46364
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_198
timestamp 1636140361
transform 1 0 55065 0 1 46363
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_199
timestamp 1636140361
transform 1 0 55062 0 1 45814
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_199
timestamp 1636140361
transform 1 0 55065 0 1 45813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_200
timestamp 1636140361
transform 1 0 55062 0 1 45574
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_200
timestamp 1636140361
transform 1 0 55065 0 1 45573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_201
timestamp 1636140361
transform 1 0 55062 0 1 45024
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_201
timestamp 1636140361
transform 1 0 55065 0 1 45023
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_202
timestamp 1636140361
transform 1 0 55062 0 1 44784
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_202
timestamp 1636140361
transform 1 0 55065 0 1 44783
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_203
timestamp 1636140361
transform 1 0 55062 0 1 44234
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_203
timestamp 1636140361
transform 1 0 55065 0 1 44233
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_204
timestamp 1636140361
transform 1 0 55062 0 1 43994
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_204
timestamp 1636140361
transform 1 0 55065 0 1 43993
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_205
timestamp 1636140361
transform 1 0 55062 0 1 43444
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_205
timestamp 1636140361
transform 1 0 55065 0 1 43443
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_206
timestamp 1636140361
transform 1 0 55062 0 1 43204
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_206
timestamp 1636140361
transform 1 0 55065 0 1 43203
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_207
timestamp 1636140361
transform 1 0 55062 0 1 42654
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_207
timestamp 1636140361
transform 1 0 55065 0 1 42653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_208
timestamp 1636140361
transform 1 0 55062 0 1 42414
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_208
timestamp 1636140361
transform 1 0 55065 0 1 42413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_209
timestamp 1636140361
transform 1 0 55062 0 1 41864
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_209
timestamp 1636140361
transform 1 0 55065 0 1 41863
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_210
timestamp 1636140361
transform 1 0 55062 0 1 41624
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_210
timestamp 1636140361
transform 1 0 55065 0 1 41623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_211
timestamp 1636140361
transform 1 0 55062 0 1 41074
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_211
timestamp 1636140361
transform 1 0 55065 0 1 41073
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_212
timestamp 1636140361
transform 1 0 55062 0 1 40834
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_212
timestamp 1636140361
transform 1 0 55065 0 1 40833
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_213
timestamp 1636140361
transform 1 0 55062 0 1 40284
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_213
timestamp 1636140361
transform 1 0 55065 0 1 40283
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_214
timestamp 1636140361
transform 1 0 55062 0 1 40044
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_214
timestamp 1636140361
transform 1 0 55065 0 1 40043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_215
timestamp 1636140361
transform 1 0 55062 0 1 39494
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_215
timestamp 1636140361
transform 1 0 55065 0 1 39493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_216
timestamp 1636140361
transform 1 0 55062 0 1 39254
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_216
timestamp 1636140361
transform 1 0 55065 0 1 39253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_217
timestamp 1636140361
transform 1 0 55062 0 1 38704
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_217
timestamp 1636140361
transform 1 0 55065 0 1 38703
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_218
timestamp 1636140361
transform 1 0 55062 0 1 38464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_218
timestamp 1636140361
transform 1 0 55065 0 1 38463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_219
timestamp 1636140361
transform 1 0 55062 0 1 37914
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_219
timestamp 1636140361
transform 1 0 55065 0 1 37913
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_220
timestamp 1636140361
transform 1 0 55062 0 1 37674
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_220
timestamp 1636140361
transform 1 0 55065 0 1 37673
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_221
timestamp 1636140361
transform 1 0 55062 0 1 37124
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_221
timestamp 1636140361
transform 1 0 55065 0 1 37123
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_222
timestamp 1636140361
transform 1 0 55062 0 1 36884
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_222
timestamp 1636140361
transform 1 0 55065 0 1 36883
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_223
timestamp 1636140361
transform 1 0 55062 0 1 36334
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_223
timestamp 1636140361
transform 1 0 55065 0 1 36333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_224
timestamp 1636140361
transform 1 0 55062 0 1 36094
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_224
timestamp 1636140361
transform 1 0 55065 0 1 36093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_225
timestamp 1636140361
transform 1 0 55062 0 1 35544
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_225
timestamp 1636140361
transform 1 0 55065 0 1 35543
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_226
timestamp 1636140361
transform 1 0 55062 0 1 35304
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_226
timestamp 1636140361
transform 1 0 55065 0 1 35303
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_227
timestamp 1636140361
transform 1 0 55062 0 1 34754
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_227
timestamp 1636140361
transform 1 0 55065 0 1 34753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_228
timestamp 1636140361
transform 1 0 55062 0 1 34514
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_228
timestamp 1636140361
transform 1 0 55065 0 1 34513
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_229
timestamp 1636140361
transform 1 0 55062 0 1 33964
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_229
timestamp 1636140361
transform 1 0 55065 0 1 33963
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_230
timestamp 1636140361
transform 1 0 55062 0 1 33724
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_230
timestamp 1636140361
transform 1 0 55065 0 1 33723
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_231
timestamp 1636140361
transform 1 0 55062 0 1 50314
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_231
timestamp 1636140361
transform 1 0 55065 0 1 50313
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_232
timestamp 1636140361
transform 1 0 55062 0 1 49764
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_232
timestamp 1636140361
transform 1 0 55065 0 1 49763
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_233
timestamp 1636140361
transform 1 0 55062 0 1 49524
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_233
timestamp 1636140361
transform 1 0 55065 0 1 49523
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_234
timestamp 1636140361
transform 1 0 55062 0 1 48974
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_234
timestamp 1636140361
transform 1 0 55065 0 1 48973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_235
timestamp 1636140361
transform 1 0 55062 0 1 48734
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_235
timestamp 1636140361
transform 1 0 55065 0 1 48733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_236
timestamp 1636140361
transform 1 0 55062 0 1 48184
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_13
timestamp 1636140361
transform 1 0 60336 0 1 63240
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_237
timestamp 1636140361
transform 1 0 60337 0 1 63245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_236
timestamp 1636140361
transform 1 0 60340 0 1 63244
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_14
timestamp 1636140361
transform 1 0 60336 0 1 66068
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_238
timestamp 1636140361
transform 1 0 60337 0 1 66073
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_237
timestamp 1636140361
transform 1 0 60340 0 1 66072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_15
timestamp 1636140361
transform 1 0 60336 0 1 64654
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_239
timestamp 1636140361
transform 1 0 60337 0 1 64659
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_238
timestamp 1636140361
transform 1 0 60340 0 1 64658
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_16
timestamp 1636140361
transform 1 0 55258 0 1 64997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_17
timestamp 1636140361
transform 1 0 55382 0 1 62470
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_18
timestamp 1636140361
transform 1 0 59332 0 1 64281
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_19
timestamp 1636140361
transform 1 0 59937 0 1 65361
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_240
timestamp 1636140361
transform 1 0 59938 0 1 65366
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_239
timestamp 1636140361
transform 1 0 59941 0 1 65365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_20
timestamp 1636140361
transform 1 0 59332 0 1 65361
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_21
timestamp 1636140361
transform 1 0 59196 0 1 64157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_22
timestamp 1636140361
transform 1 0 59937 0 1 63947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_241
timestamp 1636140361
transform 1 0 59938 0 1 63952
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_240
timestamp 1636140361
transform 1 0 59941 0 1 63951
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_23
timestamp 1636140361
transform 1 0 59196 0 1 63947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_242
timestamp 1636140361
transform 1 0 55062 0 1 60824
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_241
timestamp 1636140361
transform 1 0 55065 0 1 60823
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_243
timestamp 1636140361
transform 1 0 55062 0 1 60584
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_242
timestamp 1636140361
transform 1 0 55065 0 1 60583
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_244
timestamp 1636140361
transform 1 0 55062 0 1 60034
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_243
timestamp 1636140361
transform 1 0 55065 0 1 60033
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_245
timestamp 1636140361
transform 1 0 55062 0 1 59794
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_244
timestamp 1636140361
transform 1 0 55065 0 1 59793
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_246
timestamp 1636140361
transform 1 0 55062 0 1 59244
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_245
timestamp 1636140361
transform 1 0 55065 0 1 59243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_247
timestamp 1636140361
transform 1 0 55062 0 1 59004
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_246
timestamp 1636140361
transform 1 0 55065 0 1 59003
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_248
timestamp 1636140361
transform 1 0 55062 0 1 58454
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_247
timestamp 1636140361
transform 1 0 55065 0 1 58453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_249
timestamp 1636140361
transform 1 0 55062 0 1 58214
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_248
timestamp 1636140361
transform 1 0 55065 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_250
timestamp 1636140361
transform 1 0 55062 0 1 57664
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_249
timestamp 1636140361
transform 1 0 55065 0 1 57663
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_251
timestamp 1636140361
transform 1 0 55062 0 1 57424
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_250
timestamp 1636140361
transform 1 0 55065 0 1 57423
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_252
timestamp 1636140361
transform 1 0 55062 0 1 56874
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_251
timestamp 1636140361
transform 1 0 55065 0 1 56873
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_253
timestamp 1636140361
transform 1 0 55062 0 1 56634
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_252
timestamp 1636140361
transform 1 0 55065 0 1 56633
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_254
timestamp 1636140361
transform 1 0 55062 0 1 56084
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_253
timestamp 1636140361
transform 1 0 55065 0 1 56083
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_255
timestamp 1636140361
transform 1 0 55062 0 1 55844
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_254
timestamp 1636140361
transform 1 0 55065 0 1 55843
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_256
timestamp 1636140361
transform 1 0 55062 0 1 55294
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_255
timestamp 1636140361
transform 1 0 55065 0 1 55293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_257
timestamp 1636140361
transform 1 0 55062 0 1 55054
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_256
timestamp 1636140361
transform 1 0 55065 0 1 55053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_258
timestamp 1636140361
transform 1 0 55062 0 1 54504
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_257
timestamp 1636140361
transform 1 0 55065 0 1 54503
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_259
timestamp 1636140361
transform 1 0 55062 0 1 54264
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_258
timestamp 1636140361
transform 1 0 55065 0 1 54263
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_260
timestamp 1636140361
transform 1 0 55062 0 1 53714
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_259
timestamp 1636140361
transform 1 0 55065 0 1 53713
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_261
timestamp 1636140361
transform 1 0 55062 0 1 53474
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_260
timestamp 1636140361
transform 1 0 55065 0 1 53473
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_262
timestamp 1636140361
transform 1 0 55062 0 1 52924
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_261
timestamp 1636140361
transform 1 0 55065 0 1 52923
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_263
timestamp 1636140361
transform 1 0 55062 0 1 52684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_262
timestamp 1636140361
transform 1 0 55065 0 1 52683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_264
timestamp 1636140361
transform 1 0 55062 0 1 52134
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_263
timestamp 1636140361
transform 1 0 55065 0 1 52133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_265
timestamp 1636140361
transform 1 0 55062 0 1 51894
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_264
timestamp 1636140361
transform 1 0 55065 0 1 51893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_266
timestamp 1636140361
transform 1 0 55062 0 1 51344
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_265
timestamp 1636140361
transform 1 0 55065 0 1 51343
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_267
timestamp 1636140361
transform 1 0 55062 0 1 51104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_266
timestamp 1636140361
transform 1 0 55065 0 1 51103
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_268
timestamp 1636140361
transform 1 0 55062 0 1 50554
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_267
timestamp 1636140361
transform 1 0 55065 0 1 50553
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_24
timestamp 1636140361
transform 1 0 53640 0 1 62619
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_269
timestamp 1636140361
transform 1 0 53641 0 1 62624
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf  sky130_sram_1kbyte_1rw1r_32x256_8_pinvbuf_1
timestamp 1636140361
transform -1 0 61137 0 -1 66122
box -36 0 1536 2862
use sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0  sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0_0
timestamp 1636140361
transform -1 0 67250 0 1 10176
box 0 -60 12011 51050
use sky130_sram_1kbyte_1rw1r_32x256_8_port_address  sky130_sram_1kbyte_1rw1r_32x256_8_port_address_0
timestamp 1636140361
transform 1 0 0 0 1 10176
box 0 -490 12011 50620
use sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0  sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0_0
timestamp 1636140361
transform 1 0 12283 0 1 61526
box 0 238 41934 5702
use sky130_sram_1kbyte_1rw1r_32x256_8_port_data  sky130_sram_1kbyte_1rw1r_32x256_8_port_data_0
timestamp 1636140361
transform 1 0 12283 0 -1 9386
box -49 238 41359 9386
use sky130_sram_1kbyte_1rw1r_32x256_8_replica_bitcell_array  sky130_sram_1kbyte_1rw1r_32x256_8_replica_bitcell_array_0
timestamp 1636140361
transform 1 0 12283 0 1 9386
box -49 0 42733 52140
<< labels >>
rlabel metal3 s 53673 62626 67334 62686 4 rbl_bl_1_1
port 1 nsew
rlabel metal3 s 60702 59093 60800 59191 4 vdd
port 2 nsew
rlabel metal3 s 60702 59525 60800 59623 4 vdd
port 2 nsew
rlabel metal3 s 60320 64642 60418 64740 4 vdd
port 2 nsew
rlabel metal3 s 60270 60315 60368 60413 4 vdd
port 2 nsew
rlabel metal3 s 60270 59093 60368 59191 4 vdd
port 2 nsew
rlabel metal3 s 59492 59897 59590 59995 4 vdd
port 2 nsew
rlabel metal3 s 59492 58712 59590 58810 4 vdd
port 2 nsew
rlabel metal3 s 60702 60315 60800 60413 4 vdd
port 2 nsew
rlabel metal3 s 59492 59502 59590 59600 4 vdd
port 2 nsew
rlabel metal3 s 60270 59883 60368 59981 4 vdd
port 2 nsew
rlabel metal3 s 59467 60878 59565 60976 4 vdd
port 2 nsew
rlabel metal3 s 59492 60292 59590 60390 4 vdd
port 2 nsew
rlabel metal3 s 58635 60872 58733 60970 4 vdd
port 2 nsew
rlabel metal3 s 59492 59107 59590 59205 4 vdd
port 2 nsew
rlabel metal3 s 60702 58735 60800 58833 4 vdd
port 2 nsew
rlabel metal3 s 60702 59883 60800 59981 4 vdd
port 2 nsew
rlabel metal3 s 60270 58735 60368 58833 4 vdd
port 2 nsew
rlabel metal3 s 60270 59525 60368 59623 4 vdd
port 2 nsew
rlabel metal3 s 59888 60292 59986 60390 4 gnd
port 3 nsew
rlabel metal3 s 59888 59107 59986 59205 4 gnd
port 3 nsew
rlabel metal3 s 59888 59502 59986 59600 4 gnd
port 3 nsew
rlabel metal3 s 61127 58735 61225 58833 4 gnd
port 3 nsew
rlabel metal3 s 59888 58712 59986 58810 4 gnd
port 3 nsew
rlabel metal3 s 61127 59151 61225 59249 4 gnd
port 3 nsew
rlabel metal3 s 61127 60315 61225 60413 4 gnd
port 3 nsew
rlabel metal3 s 61127 59941 61225 60039 4 gnd
port 3 nsew
rlabel metal3 s 60320 66056 60418 66154 4 gnd
port 3 nsew
rlabel metal3 s 59888 59897 59986 59995 4 gnd
port 3 nsew
rlabel metal3 s 61127 59525 61225 59623 4 gnd
port 3 nsew
rlabel metal3 s 60320 63228 60418 63326 4 gnd
port 3 nsew
rlabel metal3 s 51360 61248 51458 61346 4 vdd
port 2 nsew
rlabel metal3 s 51429 66749 51527 66847 4 vdd
port 2 nsew
rlabel metal3 s 51417 65911 51515 66009 4 vdd
port 2 nsew
rlabel metal3 s 49993 61839 50091 61937 4 vdd
port 2 nsew
rlabel metal3 s 53351 61839 53449 61937 4 vdd
port 2 nsew
rlabel metal3 s 50112 61248 50210 61346 4 vdd
port 2 nsew
rlabel metal3 s 52489 61839 52587 61937 4 vdd
port 2 nsew
rlabel metal3 s 55944 60884 56042 60982 4 vdd
port 2 nsew
rlabel metal3 s 53737 61839 53835 61937 4 vdd
port 2 nsew
rlabel metal3 s 51984 61248 52082 61346 4 vdd
port 2 nsew
rlabel metal3 s 54552 59897 54650 59995 4 gnd
port 3 nsew
rlabel metal3 s 51429 67071 51527 67169 4 gnd
port 3 nsew
rlabel metal3 s 52103 61839 52201 61937 4 vdd
port 2 nsew
rlabel metal3 s 50736 61248 50834 61346 4 vdd
port 2 nsew
rlabel metal3 s 50181 66749 50279 66847 4 vdd
port 2 nsew
rlabel metal3 s 53232 61248 53330 61346 4 vdd
port 2 nsew
rlabel metal3 s 50251 65137 50349 65235 4 gnd
port 3 nsew
rlabel metal3 s 54552 59344 54650 59442 4 gnd
port 3 nsew
rlabel metal3 s 54552 59660 54650 59758 4 gnd
port 3 nsew
rlabel metal3 s 52920 63388 53018 63486 4 gnd
port 3 nsew
rlabel metal3 s 50169 65911 50267 66009 4 vdd
port 2 nsew
rlabel metal3 s 50855 61839 50953 61937 4 vdd
port 2 nsew
rlabel metal3 s 51499 65137 51597 65235 4 gnd
port 3 nsew
rlabel metal3 s 54552 60687 54650 60785 4 gnd
port 3 nsew
rlabel metal3 s 52747 65137 52845 65235 4 gnd
port 3 nsew
rlabel metal3 s 52665 65911 52763 66009 4 vdd
port 2 nsew
rlabel metal3 s 53856 61248 53954 61346 4 vdd
port 2 nsew
rlabel metal3 s 54552 60134 54650 60232 4 gnd
port 3 nsew
rlabel metal3 s 52677 67071 52775 67169 4 gnd
port 3 nsew
rlabel metal3 s 52677 66749 52775 66847 4 vdd
port 2 nsew
rlabel metal3 s 54552 58870 54650 58968 4 gnd
port 3 nsew
rlabel metal3 s 51241 61839 51339 61937 4 vdd
port 2 nsew
rlabel metal3 s 50424 63388 50522 63486 4 gnd
port 3 nsew
rlabel metal3 s 50181 67071 50279 67169 4 gnd
port 3 nsew
rlabel metal3 s 54918 61034 55016 61132 4 gnd
port 3 nsew
rlabel metal3 s 54552 60450 54650 60548 4 gnd
port 3 nsew
rlabel metal3 s 54552 59107 54650 59205 4 gnd
port 3 nsew
rlabel metal3 s 51672 63388 51770 63486 4 gnd
port 3 nsew
rlabel metal3 s 52608 61248 52706 61346 4 vdd
port 2 nsew
rlabel metal3 s 54552 51207 54650 51305 4 gnd
port 3 nsew
rlabel metal3 s 54552 53577 54650 53675 4 gnd
port 3 nsew
rlabel metal3 s 54552 55947 54650 56045 4 gnd
port 3 nsew
rlabel metal3 s 54552 56500 54650 56598 4 gnd
port 3 nsew
rlabel metal3 s 54552 54130 54650 54228 4 gnd
port 3 nsew
rlabel metal3 s 54552 55710 54650 55808 4 gnd
port 3 nsew
rlabel metal3 s 54552 51444 54650 51542 4 gnd
port 3 nsew
rlabel metal3 s 54552 58317 54650 58415 4 gnd
port 3 nsew
rlabel metal3 s 54552 51997 54650 52095 4 gnd
port 3 nsew
rlabel metal3 s 54552 53340 54650 53438 4 gnd
port 3 nsew
rlabel metal3 s 54552 50654 54650 50752 4 gnd
port 3 nsew
rlabel metal3 s 54552 57527 54650 57625 4 gnd
port 3 nsew
rlabel metal3 s 54552 56184 54650 56282 4 gnd
port 3 nsew
rlabel metal3 s 54552 58554 54650 58652 4 gnd
port 3 nsew
rlabel metal3 s 54552 56974 54650 57072 4 gnd
port 3 nsew
rlabel metal3 s 54552 55394 54650 55492 4 gnd
port 3 nsew
rlabel metal3 s 54552 52787 54650 52885 4 gnd
port 3 nsew
rlabel metal3 s 54552 55157 54650 55255 4 gnd
port 3 nsew
rlabel metal3 s 54552 52550 54650 52648 4 gnd
port 3 nsew
rlabel metal3 s 54552 53024 54650 53122 4 gnd
port 3 nsew
rlabel metal3 s 54552 54367 54650 54465 4 gnd
port 3 nsew
rlabel metal3 s 54552 53814 54650 53912 4 gnd
port 3 nsew
rlabel metal3 s 54552 56737 54650 56835 4 gnd
port 3 nsew
rlabel metal3 s 54552 50417 54650 50515 4 gnd
port 3 nsew
rlabel metal3 s 54552 57764 54650 57862 4 gnd
port 3 nsew
rlabel metal3 s 54552 54920 54650 55018 4 gnd
port 3 nsew
rlabel metal3 s 54552 52234 54650 52332 4 gnd
port 3 nsew
rlabel metal3 s 54552 51760 54650 51858 4 gnd
port 3 nsew
rlabel metal3 s 54552 58080 54650 58178 4 gnd
port 3 nsew
rlabel metal3 s 54552 50970 54650 51068 4 gnd
port 3 nsew
rlabel metal3 s 54552 54604 54650 54702 4 gnd
port 3 nsew
rlabel metal3 s 54552 57290 54650 57388 4 gnd
port 3 nsew
rlabel metal3 s 60270 57155 60368 57253 4 vdd
port 2 nsew
rlabel metal3 s 61127 54785 61225 54883 4 gnd
port 3 nsew
rlabel metal3 s 60702 56365 60800 56463 4 vdd
port 2 nsew
rlabel metal3 s 60270 55933 60368 56031 4 vdd
port 2 nsew
rlabel metal3 s 59888 56737 59986 56835 4 gnd
port 3 nsew
rlabel metal3 s 60270 58303 60368 58401 4 vdd
port 2 nsew
rlabel metal3 s 61127 57571 61225 57669 4 gnd
port 3 nsew
rlabel metal3 s 59492 57922 59590 58020 4 vdd
port 2 nsew
rlabel metal3 s 60270 57945 60368 58043 4 vdd
port 2 nsew
rlabel metal3 s 59888 54762 59986 54860 4 gnd
port 3 nsew
rlabel metal3 s 60702 58303 60800 58401 4 vdd
port 2 nsew
rlabel metal3 s 61127 55575 61225 55673 4 gnd
port 3 nsew
rlabel metal3 s 59888 58317 59986 58415 4 gnd
port 3 nsew
rlabel metal3 s 59888 57527 59986 57625 4 gnd
port 3 nsew
rlabel metal3 s 61127 55201 61225 55299 4 gnd
port 3 nsew
rlabel metal3 s 59492 55552 59590 55650 4 vdd
port 2 nsew
rlabel metal3 s 60702 57945 60800 58043 4 vdd
port 2 nsew
rlabel metal3 s 60702 55933 60800 56031 4 vdd
port 2 nsew
rlabel metal3 s 60702 57155 60800 57253 4 vdd
port 2 nsew
rlabel metal3 s 60270 57513 60368 57611 4 vdd
port 2 nsew
rlabel metal3 s 61127 57155 61225 57253 4 gnd
port 3 nsew
rlabel metal3 s 59888 57132 59986 57230 4 gnd
port 3 nsew
rlabel metal3 s 61127 55991 61225 56089 4 gnd
port 3 nsew
rlabel metal3 s 59492 58317 59590 58415 4 vdd
port 2 nsew
rlabel metal3 s 60702 57513 60800 57611 4 vdd
port 2 nsew
rlabel metal3 s 61127 58361 61225 58459 4 gnd
port 3 nsew
rlabel metal3 s 59888 55947 59986 56045 4 gnd
port 3 nsew
rlabel metal3 s 60702 55143 60800 55241 4 vdd
port 2 nsew
rlabel metal3 s 59492 57527 59590 57625 4 vdd
port 2 nsew
rlabel metal3 s 59888 56342 59986 56440 4 gnd
port 3 nsew
rlabel metal3 s 59492 56342 59590 56440 4 vdd
port 2 nsew
rlabel metal3 s 61127 56781 61225 56879 4 gnd
port 3 nsew
rlabel metal3 s 61127 57945 61225 58043 4 gnd
port 3 nsew
rlabel metal3 s 60270 56365 60368 56463 4 vdd
port 2 nsew
rlabel metal3 s 59888 55552 59986 55650 4 gnd
port 3 nsew
rlabel metal3 s 61127 56365 61225 56463 4 gnd
port 3 nsew
rlabel metal3 s 59888 55157 59986 55255 4 gnd
port 3 nsew
rlabel metal3 s 60270 54785 60368 54883 4 vdd
port 2 nsew
rlabel metal3 s 59492 55947 59590 56045 4 vdd
port 2 nsew
rlabel metal3 s 59492 56737 59590 56835 4 vdd
port 2 nsew
rlabel metal3 s 60270 55575 60368 55673 4 vdd
port 2 nsew
rlabel metal3 s 59492 55157 59590 55255 4 vdd
port 2 nsew
rlabel metal3 s 59888 57922 59986 58020 4 gnd
port 3 nsew
rlabel metal3 s 60702 55575 60800 55673 4 vdd
port 2 nsew
rlabel metal3 s 59492 54762 59590 54860 4 vdd
port 2 nsew
rlabel metal3 s 60270 56723 60368 56821 4 vdd
port 2 nsew
rlabel metal3 s 60270 55143 60368 55241 4 vdd
port 2 nsew
rlabel metal3 s 60702 56723 60800 56821 4 vdd
port 2 nsew
rlabel metal3 s 60702 54785 60800 54883 4 vdd
port 2 nsew
rlabel metal3 s 59492 57132 59590 57230 4 vdd
port 2 nsew
rlabel metal3 s 61127 51625 61225 51723 4 gnd
port 3 nsew
rlabel metal3 s 59492 52392 59590 52490 4 vdd
port 2 nsew
rlabel metal3 s 60702 50403 60800 50501 4 vdd
port 2 nsew
rlabel metal3 s 59492 50812 59590 50910 4 vdd
port 2 nsew
rlabel metal3 s 59492 54367 59590 54465 4 vdd
port 2 nsew
rlabel metal3 s 60270 53995 60368 54093 4 vdd
port 2 nsew
rlabel metal3 s 59492 53577 59590 53675 4 vdd
port 2 nsew
rlabel metal3 s 61127 54411 61225 54509 4 gnd
port 3 nsew
rlabel metal3 s 59888 52392 59986 52490 4 gnd
port 3 nsew
rlabel metal3 s 60270 54353 60368 54451 4 vdd
port 2 nsew
rlabel metal3 s 60270 52415 60368 52513 4 vdd
port 2 nsew
rlabel metal3 s 59888 50812 59986 50910 4 gnd
port 3 nsew
rlabel metal3 s 60702 53995 60800 54093 4 vdd
port 2 nsew
rlabel metal3 s 59492 51602 59590 51700 4 vdd
port 2 nsew
rlabel metal3 s 61127 50461 61225 50559 4 gnd
port 3 nsew
rlabel metal3 s 60702 51983 60800 52081 4 vdd
port 2 nsew
rlabel metal3 s 59492 50417 59590 50515 4 vdd
port 2 nsew
rlabel metal3 s 61127 52415 61225 52513 4 gnd
port 3 nsew
rlabel metal3 s 61127 52831 61225 52929 4 gnd
port 3 nsew
rlabel metal3 s 60702 51193 60800 51291 4 vdd
port 2 nsew
rlabel metal3 s 60702 50835 60800 50933 4 vdd
port 2 nsew
rlabel metal3 s 60270 53205 60368 53303 4 vdd
port 2 nsew
rlabel metal3 s 59888 51997 59986 52095 4 gnd
port 3 nsew
rlabel metal3 s 60270 50403 60368 50501 4 vdd
port 2 nsew
rlabel metal3 s 60702 53563 60800 53661 4 vdd
port 2 nsew
rlabel metal3 s 60702 51625 60800 51723 4 vdd
port 2 nsew
rlabel metal3 s 59888 52787 59986 52885 4 gnd
port 3 nsew
rlabel metal3 s 61127 53205 61225 53303 4 gnd
port 3 nsew
rlabel metal3 s 59888 50417 59986 50515 4 gnd
port 3 nsew
rlabel metal3 s 59888 51602 59986 51700 4 gnd
port 3 nsew
rlabel metal3 s 60702 54353 60800 54451 4 vdd
port 2 nsew
rlabel metal3 s 59492 51997 59590 52095 4 vdd
port 2 nsew
rlabel metal3 s 61127 50835 61225 50933 4 gnd
port 3 nsew
rlabel metal3 s 59492 53972 59590 54070 4 vdd
port 2 nsew
rlabel metal3 s 59888 54367 59986 54465 4 gnd
port 3 nsew
rlabel metal3 s 60702 52773 60800 52871 4 vdd
port 2 nsew
rlabel metal3 s 59888 53972 59986 54070 4 gnd
port 3 nsew
rlabel metal3 s 60270 51625 60368 51723 4 vdd
port 2 nsew
rlabel metal3 s 59492 51207 59590 51305 4 vdd
port 2 nsew
rlabel metal3 s 60702 52415 60800 52513 4 vdd
port 2 nsew
rlabel metal3 s 59888 51207 59986 51305 4 gnd
port 3 nsew
rlabel metal3 s 61127 51251 61225 51349 4 gnd
port 3 nsew
rlabel metal3 s 59888 53577 59986 53675 4 gnd
port 3 nsew
rlabel metal3 s 60270 51193 60368 51291 4 vdd
port 2 nsew
rlabel metal3 s 60702 53205 60800 53303 4 vdd
port 2 nsew
rlabel metal3 s 59888 53182 59986 53280 4 gnd
port 3 nsew
rlabel metal3 s 60270 51983 60368 52081 4 vdd
port 2 nsew
rlabel metal3 s 61127 53995 61225 54093 4 gnd
port 3 nsew
rlabel metal3 s 60270 53563 60368 53661 4 vdd
port 2 nsew
rlabel metal3 s 59492 52787 59590 52885 4 vdd
port 2 nsew
rlabel metal3 s 61127 52041 61225 52139 4 gnd
port 3 nsew
rlabel metal3 s 61127 53621 61225 53719 4 gnd
port 3 nsew
rlabel metal3 s 60270 50835 60368 50933 4 vdd
port 2 nsew
rlabel metal3 s 60270 52773 60368 52871 4 vdd
port 2 nsew
rlabel metal3 s 59492 53182 59590 53280 4 vdd
port 2 nsew
rlabel metal3 s 43367 61839 43465 61937 4 vdd
port 2 nsew
rlabel metal3 s 44615 61839 44713 61937 4 vdd
port 2 nsew
rlabel metal3 s 47673 65911 47771 66009 4 vdd
port 2 nsew
rlabel metal3 s 49607 61839 49705 61937 4 vdd
port 2 nsew
rlabel metal3 s 42000 61248 42098 61346 4 vdd
port 2 nsew
rlabel metal3 s 46437 66749 46535 66847 4 vdd
port 2 nsew
rlabel metal3 s 44011 65137 44109 65235 4 gnd
port 3 nsew
rlabel metal3 s 48745 61839 48843 61937 4 vdd
port 2 nsew
rlabel metal3 s 49176 63388 49274 63486 4 gnd
port 3 nsew
rlabel metal3 s 46249 61839 46347 61937 4 vdd
port 2 nsew
rlabel metal3 s 44496 61248 44594 61346 4 vdd
port 2 nsew
rlabel metal3 s 42505 61839 42603 61937 4 vdd
port 2 nsew
rlabel metal3 s 48864 61248 48962 61346 4 vdd
port 2 nsew
rlabel metal3 s 48240 61248 48338 61346 4 vdd
port 2 nsew
rlabel metal3 s 49003 65137 49101 65235 4 gnd
port 3 nsew
rlabel metal3 s 43753 61839 43851 61937 4 vdd
port 2 nsew
rlabel metal3 s 42119 61839 42217 61937 4 vdd
port 2 nsew
rlabel metal3 s 43929 65911 44027 66009 4 vdd
port 2 nsew
rlabel metal3 s 46425 65911 46523 66009 4 vdd
port 2 nsew
rlabel metal3 s 42693 67071 42791 67169 4 gnd
port 3 nsew
rlabel metal3 s 45120 61248 45218 61346 4 vdd
port 2 nsew
rlabel metal3 s 47928 63388 48026 63486 4 gnd
port 3 nsew
rlabel metal3 s 45259 65137 45357 65235 4 gnd
port 3 nsew
rlabel metal3 s 44184 63388 44282 63486 4 gnd
port 3 nsew
rlabel metal3 s 46992 61248 47090 61346 4 vdd
port 2 nsew
rlabel metal3 s 47497 61839 47595 61937 4 vdd
port 2 nsew
rlabel metal3 s 45001 61839 45099 61937 4 vdd
port 2 nsew
rlabel metal3 s 45189 67071 45287 67169 4 gnd
port 3 nsew
rlabel metal3 s 42763 65137 42861 65235 4 gnd
port 3 nsew
rlabel metal3 s 43872 61248 43970 61346 4 vdd
port 2 nsew
rlabel metal3 s 43941 67071 44039 67169 4 gnd
port 3 nsew
rlabel metal3 s 47111 61839 47209 61937 4 vdd
port 2 nsew
rlabel metal3 s 45189 66749 45287 66847 4 vdd
port 2 nsew
rlabel metal3 s 46368 61248 46466 61346 4 vdd
port 2 nsew
rlabel metal3 s 48933 66749 49031 66847 4 vdd
port 2 nsew
rlabel metal3 s 45177 65911 45275 66009 4 vdd
port 2 nsew
rlabel metal3 s 45744 61248 45842 61346 4 vdd
port 2 nsew
rlabel metal3 s 47685 67071 47783 67169 4 gnd
port 3 nsew
rlabel metal3 s 42624 61248 42722 61346 4 vdd
port 2 nsew
rlabel metal3 s 49488 61248 49586 61346 4 vdd
port 2 nsew
rlabel metal3 s 42681 65911 42779 66009 4 vdd
port 2 nsew
rlabel metal3 s 47616 61248 47714 61346 4 vdd
port 2 nsew
rlabel metal3 s 43941 66749 44039 66847 4 vdd
port 2 nsew
rlabel metal3 s 48933 67071 49031 67169 4 gnd
port 3 nsew
rlabel metal3 s 42693 66749 42791 66847 4 vdd
port 2 nsew
rlabel metal3 s 46680 63388 46778 63486 4 gnd
port 3 nsew
rlabel metal3 s 48359 61839 48457 61937 4 vdd
port 2 nsew
rlabel metal3 s 46437 67071 46535 67169 4 gnd
port 3 nsew
rlabel metal3 s 45432 63388 45530 63486 4 gnd
port 3 nsew
rlabel metal3 s 41688 63388 41786 63486 4 gnd
port 3 nsew
rlabel metal3 s 46507 65137 46605 65235 4 gnd
port 3 nsew
rlabel metal3 s 42936 63388 43034 63486 4 gnd
port 3 nsew
rlabel metal3 s 45863 61839 45961 61937 4 vdd
port 2 nsew
rlabel metal3 s 43248 61248 43346 61346 4 vdd
port 2 nsew
rlabel metal3 s 48921 65911 49019 66009 4 vdd
port 2 nsew
rlabel metal3 s 47685 66749 47783 66847 4 vdd
port 2 nsew
rlabel metal3 s 47755 65137 47853 65235 4 gnd
port 3 nsew
rlabel metal3 s 40267 65137 40365 65235 4 gnd
port 3 nsew
rlabel metal3 s 41376 61248 41474 61346 4 vdd
port 2 nsew
rlabel metal3 s 41257 61839 41355 61937 4 vdd
port 2 nsew
rlabel metal3 s 36265 61839 36363 61937 4 vdd
port 2 nsew
rlabel metal3 s 35017 61839 35115 61937 4 vdd
port 2 nsew
rlabel metal3 s 39192 63388 39290 63486 4 gnd
port 3 nsew
rlabel metal3 s 33957 66749 34055 66847 4 vdd
port 2 nsew
rlabel metal3 s 33888 61248 33986 61346 4 vdd
port 2 nsew
rlabel metal3 s 38949 66749 39047 66847 4 vdd
port 2 nsew
rlabel metal3 s 37944 63388 38042 63486 4 gnd
port 3 nsew
rlabel metal3 s 37701 66749 37799 66847 4 vdd
port 2 nsew
rlabel metal3 s 36384 61248 36482 61346 4 vdd
port 2 nsew
rlabel metal3 s 33945 65911 34043 66009 4 vdd
port 2 nsew
rlabel metal3 s 35275 65137 35373 65235 4 gnd
port 3 nsew
rlabel metal3 s 34512 61248 34610 61346 4 vdd
port 2 nsew
rlabel metal3 s 41445 67071 41543 67169 4 gnd
port 3 nsew
rlabel metal3 s 39504 61248 39602 61346 4 vdd
port 2 nsew
rlabel metal3 s 38761 61839 38859 61937 4 vdd
port 2 nsew
rlabel metal3 s 35448 63388 35546 63486 4 gnd
port 3 nsew
rlabel metal3 s 35760 61248 35858 61346 4 vdd
port 2 nsew
rlabel metal3 s 38375 61839 38473 61937 4 vdd
port 2 nsew
rlabel metal3 s 40185 65911 40283 66009 4 vdd
port 2 nsew
rlabel metal3 s 35205 67071 35303 67169 4 gnd
port 3 nsew
rlabel metal3 s 41433 65911 41531 66009 4 vdd
port 2 nsew
rlabel metal3 s 34200 63388 34298 63486 4 gnd
port 3 nsew
rlabel metal3 s 35136 61248 35234 61346 4 vdd
port 2 nsew
rlabel metal3 s 40752 61248 40850 61346 4 vdd
port 2 nsew
rlabel metal3 s 34631 61839 34729 61937 4 vdd
port 2 nsew
rlabel metal3 s 41445 66749 41543 66847 4 vdd
port 2 nsew
rlabel metal3 s 40197 66749 40295 66847 4 vdd
port 2 nsew
rlabel metal3 s 35205 66749 35303 66847 4 vdd
port 2 nsew
rlabel metal3 s 35879 61839 35977 61937 4 vdd
port 2 nsew
rlabel metal3 s 38937 65911 39035 66009 4 vdd
port 2 nsew
rlabel metal3 s 40009 61839 40107 61937 4 vdd
port 2 nsew
rlabel metal3 s 37127 61839 37225 61937 4 vdd
port 2 nsew
rlabel metal3 s 38256 61248 38354 61346 4 vdd
port 2 nsew
rlabel metal3 s 40871 61839 40969 61937 4 vdd
port 2 nsew
rlabel metal3 s 33769 61839 33867 61937 4 vdd
port 2 nsew
rlabel metal3 s 40197 67071 40295 67169 4 gnd
port 3 nsew
rlabel metal3 s 39019 65137 39117 65235 4 gnd
port 3 nsew
rlabel metal3 s 36453 66749 36551 66847 4 vdd
port 2 nsew
rlabel metal3 s 40128 61248 40226 61346 4 vdd
port 2 nsew
rlabel metal3 s 37771 65137 37869 65235 4 gnd
port 3 nsew
rlabel metal3 s 36453 67071 36551 67169 4 gnd
port 3 nsew
rlabel metal3 s 41515 65137 41613 65235 4 gnd
port 3 nsew
rlabel metal3 s 37701 67071 37799 67169 4 gnd
port 3 nsew
rlabel metal3 s 37008 61248 37106 61346 4 vdd
port 2 nsew
rlabel metal3 s 40440 63388 40538 63486 4 gnd
port 3 nsew
rlabel metal3 s 37689 65911 37787 66009 4 vdd
port 2 nsew
rlabel metal3 s 36696 63388 36794 63486 4 gnd
port 3 nsew
rlabel metal3 s 35193 65911 35291 66009 4 vdd
port 2 nsew
rlabel metal3 s 34027 65137 34125 65235 4 gnd
port 3 nsew
rlabel metal3 s 38949 67071 39047 67169 4 gnd
port 3 nsew
rlabel metal3 s 37513 61839 37611 61937 4 vdd
port 2 nsew
rlabel metal3 s 37632 61248 37730 61346 4 vdd
port 2 nsew
rlabel metal3 s 38880 61248 38978 61346 4 vdd
port 2 nsew
rlabel metal3 s 33957 67071 34055 67169 4 gnd
port 3 nsew
rlabel metal3 s 36523 65137 36621 65235 4 gnd
port 3 nsew
rlabel metal3 s 39623 61839 39721 61937 4 vdd
port 2 nsew
rlabel metal3 s 36441 65911 36539 66009 4 vdd
port 2 nsew
rlabel metal3 s 59888 50022 59986 50120 4 gnd
port 3 nsew
rlabel metal3 s 61127 48881 61225 48979 4 gnd
port 3 nsew
rlabel metal3 s 61127 47301 61225 47399 4 gnd
port 3 nsew
rlabel metal3 s 59492 47652 59590 47750 4 vdd
port 2 nsew
rlabel metal3 s 60270 46453 60368 46551 4 vdd
port 2 nsew
rlabel metal3 s 61127 46885 61225 46983 4 gnd
port 3 nsew
rlabel metal3 s 60702 50045 60800 50143 4 vdd
port 2 nsew
rlabel metal3 s 60702 48033 60800 48131 4 vdd
port 2 nsew
rlabel metal3 s 60270 46885 60368 46983 4 vdd
port 2 nsew
rlabel metal3 s 61127 48091 61225 48189 4 gnd
port 3 nsew
rlabel metal3 s 60270 47243 60368 47341 4 vdd
port 2 nsew
rlabel metal3 s 61127 48465 61225 48563 4 gnd
port 3 nsew
rlabel metal3 s 60270 48465 60368 48563 4 vdd
port 2 nsew
rlabel metal3 s 60702 49613 60800 49711 4 vdd
port 2 nsew
rlabel metal3 s 59888 48047 59986 48145 4 gnd
port 3 nsew
rlabel metal3 s 59888 46467 59986 46565 4 gnd
port 3 nsew
rlabel metal3 s 60270 47675 60368 47773 4 vdd
port 2 nsew
rlabel metal3 s 61127 47675 61225 47773 4 gnd
port 3 nsew
rlabel metal3 s 59492 47257 59590 47355 4 vdd
port 2 nsew
rlabel metal3 s 60702 47243 60800 47341 4 vdd
port 2 nsew
rlabel metal3 s 59888 48837 59986 48935 4 gnd
port 3 nsew
rlabel metal3 s 59888 47257 59986 47355 4 gnd
port 3 nsew
rlabel metal3 s 59492 48047 59590 48145 4 vdd
port 2 nsew
rlabel metal3 s 61127 49671 61225 49769 4 gnd
port 3 nsew
rlabel metal3 s 59492 50022 59590 50120 4 vdd
port 2 nsew
rlabel metal3 s 59492 46467 59590 46565 4 vdd
port 2 nsew
rlabel metal3 s 60702 48823 60800 48921 4 vdd
port 2 nsew
rlabel metal3 s 59888 48442 59986 48540 4 gnd
port 3 nsew
rlabel metal3 s 60270 48033 60368 48131 4 vdd
port 2 nsew
rlabel metal3 s 60702 47675 60800 47773 4 vdd
port 2 nsew
rlabel metal3 s 61127 46511 61225 46609 4 gnd
port 3 nsew
rlabel metal3 s 60702 48465 60800 48563 4 vdd
port 2 nsew
rlabel metal3 s 60702 49255 60800 49353 4 vdd
port 2 nsew
rlabel metal3 s 60702 46885 60800 46983 4 vdd
port 2 nsew
rlabel metal3 s 59492 48442 59590 48540 4 vdd
port 2 nsew
rlabel metal3 s 59492 49627 59590 49725 4 vdd
port 2 nsew
rlabel metal3 s 59888 49627 59986 49725 4 gnd
port 3 nsew
rlabel metal3 s 59888 49232 59986 49330 4 gnd
port 3 nsew
rlabel metal3 s 60270 50045 60368 50143 4 vdd
port 2 nsew
rlabel metal3 s 59492 48837 59590 48935 4 vdd
port 2 nsew
rlabel metal3 s 59888 47652 59986 47750 4 gnd
port 3 nsew
rlabel metal3 s 61127 49255 61225 49353 4 gnd
port 3 nsew
rlabel metal3 s 60702 46453 60800 46551 4 vdd
port 2 nsew
rlabel metal3 s 60270 49255 60368 49353 4 vdd
port 2 nsew
rlabel metal3 s 59492 46862 59590 46960 4 vdd
port 2 nsew
rlabel metal3 s 59888 46862 59986 46960 4 gnd
port 3 nsew
rlabel metal3 s 60270 49613 60368 49711 4 vdd
port 2 nsew
rlabel metal3 s 61127 50045 61225 50143 4 gnd
port 3 nsew
rlabel metal3 s 59492 49232 59590 49330 4 vdd
port 2 nsew
rlabel metal3 s 60270 48823 60368 48921 4 vdd
port 2 nsew
rlabel metal3 s 60270 46095 60368 46193 4 vdd
port 2 nsew
rlabel metal3 s 59492 43307 59590 43405 4 vdd
port 2 nsew
rlabel metal3 s 60702 44083 60800 44181 4 vdd
port 2 nsew
rlabel metal3 s 61127 42935 61225 43033 4 gnd
port 3 nsew
rlabel metal3 s 60270 42935 60368 43033 4 vdd
port 2 nsew
rlabel metal3 s 61127 44141 61225 44239 4 gnd
port 3 nsew
rlabel metal3 s 60270 43725 60368 43823 4 vdd
port 2 nsew
rlabel metal3 s 61127 45721 61225 45819 4 gnd
port 3 nsew
rlabel metal3 s 60702 42935 60800 43033 4 vdd
port 2 nsew
rlabel metal3 s 60270 43293 60368 43391 4 vdd
port 2 nsew
rlabel metal3 s 60702 42145 60800 42243 4 vdd
port 2 nsew
rlabel metal3 s 59492 44097 59590 44195 4 vdd
port 2 nsew
rlabel metal3 s 59888 44097 59986 44195 4 gnd
port 3 nsew
rlabel metal3 s 61127 45305 61225 45403 4 gnd
port 3 nsew
rlabel metal3 s 59492 44887 59590 44985 4 vdd
port 2 nsew
rlabel metal3 s 60702 46095 60800 46193 4 vdd
port 2 nsew
rlabel metal3 s 60270 42503 60368 42601 4 vdd
port 2 nsew
rlabel metal3 s 59492 42912 59590 43010 4 vdd
port 2 nsew
rlabel metal3 s 59888 42912 59986 43010 4 gnd
port 3 nsew
rlabel metal3 s 60270 45305 60368 45403 4 vdd
port 2 nsew
rlabel metal3 s 61127 46095 61225 46193 4 gnd
port 3 nsew
rlabel metal3 s 59888 43702 59986 43800 4 gnd
port 3 nsew
rlabel metal3 s 60702 42503 60800 42601 4 vdd
port 2 nsew
rlabel metal3 s 61127 42561 61225 42659 4 gnd
port 3 nsew
rlabel metal3 s 60702 45663 60800 45761 4 vdd
port 2 nsew
rlabel metal3 s 59888 45677 59986 45775 4 gnd
port 3 nsew
rlabel metal3 s 60702 43725 60800 43823 4 vdd
port 2 nsew
rlabel metal3 s 61127 43725 61225 43823 4 gnd
port 3 nsew
rlabel metal3 s 59492 45677 59590 45775 4 vdd
port 2 nsew
rlabel metal3 s 61127 43351 61225 43449 4 gnd
port 3 nsew
rlabel metal3 s 60270 44083 60368 44181 4 vdd
port 2 nsew
rlabel metal3 s 59492 44492 59590 44590 4 vdd
port 2 nsew
rlabel metal3 s 60702 44515 60800 44613 4 vdd
port 2 nsew
rlabel metal3 s 59492 42517 59590 42615 4 vdd
port 2 nsew
rlabel metal3 s 60702 43293 60800 43391 4 vdd
port 2 nsew
rlabel metal3 s 60270 45663 60368 45761 4 vdd
port 2 nsew
rlabel metal3 s 60270 42145 60368 42243 4 vdd
port 2 nsew
rlabel metal3 s 59888 44887 59986 44985 4 gnd
port 3 nsew
rlabel metal3 s 59888 42517 59986 42615 4 gnd
port 3 nsew
rlabel metal3 s 59492 42122 59590 42220 4 vdd
port 2 nsew
rlabel metal3 s 59888 43307 59986 43405 4 gnd
port 3 nsew
rlabel metal3 s 61127 42145 61225 42243 4 gnd
port 3 nsew
rlabel metal3 s 59888 45282 59986 45380 4 gnd
port 3 nsew
rlabel metal3 s 59492 43702 59590 43800 4 vdd
port 2 nsew
rlabel metal3 s 61127 44931 61225 45029 4 gnd
port 3 nsew
rlabel metal3 s 60702 45305 60800 45403 4 vdd
port 2 nsew
rlabel metal3 s 59492 45282 59590 45380 4 vdd
port 2 nsew
rlabel metal3 s 59888 42122 59986 42220 4 gnd
port 3 nsew
rlabel metal3 s 60270 44515 60368 44613 4 vdd
port 2 nsew
rlabel metal3 s 60270 44873 60368 44971 4 vdd
port 2 nsew
rlabel metal3 s 59888 44492 59986 44590 4 gnd
port 3 nsew
rlabel metal3 s 60702 44873 60800 44971 4 vdd
port 2 nsew
rlabel metal3 s 59492 46072 59590 46170 4 vdd
port 2 nsew
rlabel metal3 s 59888 46072 59986 46170 4 gnd
port 3 nsew
rlabel metal3 s 61127 44515 61225 44613 4 gnd
port 3 nsew
rlabel metal3 s 54552 41964 54650 42062 4 gnd
port 3 nsew
rlabel metal3 s 54552 43860 54650 43958 4 gnd
port 3 nsew
rlabel metal3 s 54552 45914 54650 46012 4 gnd
port 3 nsew
rlabel metal3 s 54552 44097 54650 44195 4 gnd
port 3 nsew
rlabel metal3 s 54552 43307 54650 43405 4 gnd
port 3 nsew
rlabel metal3 s 54552 49074 54650 49172 4 gnd
port 3 nsew
rlabel metal3 s 54552 46230 54650 46328 4 gnd
port 3 nsew
rlabel metal3 s 54552 49627 54650 49725 4 gnd
port 3 nsew
rlabel metal3 s 54552 45124 54650 45222 4 gnd
port 3 nsew
rlabel metal3 s 54552 43544 54650 43642 4 gnd
port 3 nsew
rlabel metal3 s 54552 47020 54650 47118 4 gnd
port 3 nsew
rlabel metal3 s 54552 42280 54650 42378 4 gnd
port 3 nsew
rlabel metal3 s 54552 49390 54650 49488 4 gnd
port 3 nsew
rlabel metal3 s 54552 47257 54650 47355 4 gnd
port 3 nsew
rlabel metal3 s 54552 48284 54650 48382 4 gnd
port 3 nsew
rlabel metal3 s 54552 45677 54650 45775 4 gnd
port 3 nsew
rlabel metal3 s 54552 46704 54650 46802 4 gnd
port 3 nsew
rlabel metal3 s 54552 42517 54650 42615 4 gnd
port 3 nsew
rlabel metal3 s 54552 47494 54650 47592 4 gnd
port 3 nsew
rlabel metal3 s 54552 44334 54650 44432 4 gnd
port 3 nsew
rlabel metal3 s 54552 48047 54650 48145 4 gnd
port 3 nsew
rlabel metal3 s 54552 48837 54650 48935 4 gnd
port 3 nsew
rlabel metal3 s 54552 48600 54650 48698 4 gnd
port 3 nsew
rlabel metal3 s 54552 45440 54650 45538 4 gnd
port 3 nsew
rlabel metal3 s 54552 43070 54650 43168 4 gnd
port 3 nsew
rlabel metal3 s 54552 50180 54650 50278 4 gnd
port 3 nsew
rlabel metal3 s 54552 47810 54650 47908 4 gnd
port 3 nsew
rlabel metal3 s 54552 46467 54650 46565 4 gnd
port 3 nsew
rlabel metal3 s 54552 42754 54650 42852 4 gnd
port 3 nsew
rlabel metal3 s 54552 44887 54650 44985 4 gnd
port 3 nsew
rlabel metal3 s 54552 49864 54650 49962 4 gnd
port 3 nsew
rlabel metal3 s 54552 44650 54650 44748 4 gnd
port 3 nsew
rlabel metal3 s 54552 35170 54650 35268 4 gnd
port 3 nsew
rlabel metal3 s 55944 35407 56042 35505 4 vdd
port 2 nsew
rlabel metal3 s 54552 41727 54650 41825 4 gnd
port 3 nsew
rlabel metal3 s 54552 37540 54650 37638 4 gnd
port 3 nsew
rlabel metal3 s 54552 35960 54650 36058 4 gnd
port 3 nsew
rlabel metal3 s 54552 39120 54650 39218 4 gnd
port 3 nsew
rlabel metal3 s 54552 41490 54650 41588 4 gnd
port 3 nsew
rlabel metal3 s 54552 36197 54650 36295 4 gnd
port 3 nsew
rlabel metal3 s 54552 35644 54650 35742 4 gnd
port 3 nsew
rlabel metal3 s 54552 39910 54650 40008 4 gnd
port 3 nsew
rlabel metal3 s 54552 36987 54650 37085 4 gnd
port 3 nsew
rlabel metal3 s 54552 34617 54650 34715 4 gnd
port 3 nsew
rlabel metal3 s 54552 34380 54650 34478 4 gnd
port 3 nsew
rlabel metal3 s 54552 38804 54650 38902 4 gnd
port 3 nsew
rlabel metal3 s 54552 37224 54650 37322 4 gnd
port 3 nsew
rlabel metal3 s 54552 34064 54650 34162 4 gnd
port 3 nsew
rlabel metal3 s 54552 38330 54650 38428 4 gnd
port 3 nsew
rlabel metal3 s 54552 35407 54650 35505 4 gnd
port 3 nsew
rlabel metal3 s 54552 40700 54650 40798 4 gnd
port 3 nsew
rlabel metal3 s 54552 34854 54650 34952 4 gnd
port 3 nsew
rlabel metal3 s 54552 39357 54650 39455 4 gnd
port 3 nsew
rlabel metal3 s 54552 33827 54650 33925 4 gnd
port 3 nsew
rlabel metal3 s 54552 39594 54650 39692 4 gnd
port 3 nsew
rlabel metal3 s 54552 36750 54650 36848 4 gnd
port 3 nsew
rlabel metal3 s 54552 38014 54650 38112 4 gnd
port 3 nsew
rlabel metal3 s 54552 38567 54650 38665 4 gnd
port 3 nsew
rlabel metal3 s 54552 40147 54650 40245 4 gnd
port 3 nsew
rlabel metal3 s 57592 35407 57690 35505 4 gnd
port 3 nsew
rlabel metal3 s 54552 37777 54650 37875 4 gnd
port 3 nsew
rlabel metal3 s 54552 33590 54650 33688 4 gnd
port 3 nsew
rlabel metal3 s 54552 36434 54650 36532 4 gnd
port 3 nsew
rlabel metal3 s 54552 40384 54650 40482 4 gnd
port 3 nsew
rlabel metal3 s 54552 41174 54650 41272 4 gnd
port 3 nsew
rlabel metal3 s 54552 40937 54650 41035 4 gnd
port 3 nsew
rlabel metal3 s 61127 41355 61225 41453 4 gnd
port 3 nsew
rlabel metal3 s 59492 39357 59590 39455 4 vdd
port 2 nsew
rlabel metal3 s 61127 38611 61225 38709 4 gnd
port 3 nsew
rlabel metal3 s 60270 37763 60368 37861 4 vdd
port 2 nsew
rlabel metal3 s 60702 38195 60800 38293 4 vdd
port 2 nsew
rlabel metal3 s 60270 39775 60368 39873 4 vdd
port 2 nsew
rlabel metal3 s 61127 41771 61225 41869 4 gnd
port 3 nsew
rlabel metal3 s 60270 40923 60368 41021 4 vdd
port 2 nsew
rlabel metal3 s 59888 37777 59986 37875 4 gnd
port 3 nsew
rlabel metal3 s 59888 41727 59986 41825 4 gnd
port 3 nsew
rlabel metal3 s 59492 38172 59590 38270 4 vdd
port 2 nsew
rlabel metal3 s 59888 41332 59986 41430 4 gnd
port 3 nsew
rlabel metal3 s 60270 38553 60368 38651 4 vdd
port 2 nsew
rlabel metal3 s 60702 41355 60800 41453 4 vdd
port 2 nsew
rlabel metal3 s 59492 40937 59590 41035 4 vdd
port 2 nsew
rlabel metal3 s 59888 38172 59986 38270 4 gnd
port 3 nsew
rlabel metal3 s 60702 39343 60800 39441 4 vdd
port 2 nsew
rlabel metal3 s 59492 41332 59590 41430 4 vdd
port 2 nsew
rlabel metal3 s 61127 40981 61225 41079 4 gnd
port 3 nsew
rlabel metal3 s 60702 40923 60800 41021 4 vdd
port 2 nsew
rlabel metal3 s 59492 38962 59590 39060 4 vdd
port 2 nsew
rlabel metal3 s 59492 38567 59590 38665 4 vdd
port 2 nsew
rlabel metal3 s 59888 38567 59986 38665 4 gnd
port 3 nsew
rlabel metal3 s 59888 40147 59986 40245 4 gnd
port 3 nsew
rlabel metal3 s 61127 39401 61225 39499 4 gnd
port 3 nsew
rlabel metal3 s 60270 40565 60368 40663 4 vdd
port 2 nsew
rlabel metal3 s 59492 39752 59590 39850 4 vdd
port 2 nsew
rlabel metal3 s 60702 39775 60800 39873 4 vdd
port 2 nsew
rlabel metal3 s 59888 39357 59986 39455 4 gnd
port 3 nsew
rlabel metal3 s 60270 41355 60368 41453 4 vdd
port 2 nsew
rlabel metal3 s 60702 41713 60800 41811 4 vdd
port 2 nsew
rlabel metal3 s 61127 39775 61225 39873 4 gnd
port 3 nsew
rlabel metal3 s 59492 40147 59590 40245 4 vdd
port 2 nsew
rlabel metal3 s 59492 40542 59590 40640 4 vdd
port 2 nsew
rlabel metal3 s 60270 41713 60368 41811 4 vdd
port 2 nsew
rlabel metal3 s 61127 40191 61225 40289 4 gnd
port 3 nsew
rlabel metal3 s 61127 40565 61225 40663 4 gnd
port 3 nsew
rlabel metal3 s 60702 38985 60800 39083 4 vdd
port 2 nsew
rlabel metal3 s 59492 41727 59590 41825 4 vdd
port 2 nsew
rlabel metal3 s 59888 39752 59986 39850 4 gnd
port 3 nsew
rlabel metal3 s 60702 40565 60800 40663 4 vdd
port 2 nsew
rlabel metal3 s 60270 40133 60368 40231 4 vdd
port 2 nsew
rlabel metal3 s 61127 37821 61225 37919 4 gnd
port 3 nsew
rlabel metal3 s 60702 38553 60800 38651 4 vdd
port 2 nsew
rlabel metal3 s 61127 38985 61225 39083 4 gnd
port 3 nsew
rlabel metal3 s 60270 39343 60368 39441 4 vdd
port 2 nsew
rlabel metal3 s 59888 38962 59986 39060 4 gnd
port 3 nsew
rlabel metal3 s 60702 40133 60800 40231 4 vdd
port 2 nsew
rlabel metal3 s 60702 37763 60800 37861 4 vdd
port 2 nsew
rlabel metal3 s 59888 40542 59986 40640 4 gnd
port 3 nsew
rlabel metal3 s 61127 38195 61225 38293 4 gnd
port 3 nsew
rlabel metal3 s 60270 38195 60368 38293 4 vdd
port 2 nsew
rlabel metal3 s 59888 40937 59986 41035 4 gnd
port 3 nsew
rlabel metal3 s 60270 38985 60368 39083 4 vdd
port 2 nsew
rlabel metal3 s 59492 37777 59590 37875 4 vdd
port 2 nsew
rlabel metal3 s 60702 36615 60800 36713 4 vdd
port 2 nsew
rlabel metal3 s 59492 36592 59590 36690 4 vdd
port 2 nsew
rlabel metal3 s 60702 35035 60800 35133 4 vdd
port 2 nsew
rlabel metal3 s 60270 34245 60368 34343 4 vdd
port 2 nsew
rlabel metal3 s 59888 35802 59986 35900 4 gnd
port 3 nsew
rlabel metal3 s 59492 34617 59590 34715 4 vdd
port 2 nsew
rlabel metal3 s 59888 36197 59986 36295 4 gnd
port 3 nsew
rlabel metal3 s 60702 36973 60800 37071 4 vdd
port 2 nsew
rlabel metal3 s 59888 35407 59986 35505 4 gnd
port 3 nsew
rlabel metal3 s 59888 36592 59986 36690 4 gnd
port 3 nsew
rlabel metal3 s 61127 34245 61225 34343 4 gnd
port 3 nsew
rlabel metal3 s 59492 36197 59590 36295 4 vdd
port 2 nsew
rlabel metal3 s 60270 34603 60368 34701 4 vdd
port 2 nsew
rlabel metal3 s 60270 36973 60368 37071 4 vdd
port 2 nsew
rlabel metal3 s 59888 37382 59986 37480 4 gnd
port 3 nsew
rlabel metal3 s 60702 36183 60800 36281 4 vdd
port 2 nsew
rlabel metal3 s 61127 37405 61225 37503 4 gnd
port 3 nsew
rlabel metal3 s 60270 35393 60368 35491 4 vdd
port 2 nsew
rlabel metal3 s 60702 35825 60800 35923 4 vdd
port 2 nsew
rlabel metal3 s 60702 37405 60800 37503 4 vdd
port 2 nsew
rlabel metal3 s 60270 37405 60368 37503 4 vdd
port 2 nsew
rlabel metal3 s 58635 35391 58733 35489 4 vdd
port 2 nsew
rlabel metal3 s 60702 33813 60800 33911 4 vdd
port 2 nsew
rlabel metal3 s 60702 34245 60800 34343 4 vdd
port 2 nsew
rlabel metal3 s 61127 35825 61225 35923 4 gnd
port 3 nsew
rlabel metal3 s 61127 35451 61225 35549 4 gnd
port 3 nsew
rlabel metal3 s 59492 35407 59590 35505 4 vdd
port 2 nsew
rlabel metal3 s 61127 35035 61225 35133 4 gnd
port 3 nsew
rlabel metal3 s 60270 36615 60368 36713 4 vdd
port 2 nsew
rlabel metal3 s 61127 36241 61225 36339 4 gnd
port 3 nsew
rlabel metal3 s 59888 35012 59986 35110 4 gnd
port 3 nsew
rlabel metal3 s 60270 35825 60368 35923 4 vdd
port 2 nsew
rlabel metal3 s 59492 34222 59590 34320 4 vdd
port 2 nsew
rlabel metal3 s 59888 33827 59986 33925 4 gnd
port 3 nsew
rlabel metal3 s 59492 37382 59590 37480 4 vdd
port 2 nsew
rlabel metal3 s 61127 34661 61225 34759 4 gnd
port 3 nsew
rlabel metal3 s 59492 35802 59590 35900 4 vdd
port 2 nsew
rlabel metal3 s 59888 34222 59986 34320 4 gnd
port 3 nsew
rlabel metal3 s 60270 35035 60368 35133 4 vdd
port 2 nsew
rlabel metal3 s 60270 33813 60368 33911 4 vdd
port 2 nsew
rlabel metal3 s 59492 33827 59590 33925 4 vdd
port 2 nsew
rlabel metal3 s 59888 34617 59986 34715 4 gnd
port 3 nsew
rlabel metal3 s 59492 35012 59590 35110 4 vdd
port 2 nsew
rlabel metal3 s 61127 33871 61225 33969 4 gnd
port 3 nsew
rlabel metal3 s 59492 36987 59590 37085 4 vdd
port 2 nsew
rlabel metal3 s 59888 36987 59986 37085 4 gnd
port 3 nsew
rlabel metal3 s 60702 35393 60800 35491 4 vdd
port 2 nsew
rlabel metal3 s 60702 34603 60800 34701 4 vdd
port 2 nsew
rlabel metal3 s 61127 36615 61225 36713 4 gnd
port 3 nsew
rlabel metal3 s 61127 37031 61225 37129 4 gnd
port 3 nsew
rlabel metal3 s 59060 35392 59158 35490 4 gnd
port 3 nsew
rlabel metal3 s 60270 36183 60368 36281 4 vdd
port 2 nsew
rlabel metal3 s 32135 61839 32233 61937 4 vdd
port 2 nsew
rlabel metal3 s 28953 65911 29051 66009 4 vdd
port 2 nsew
rlabel metal3 s 32779 65137 32877 65235 4 gnd
port 3 nsew
rlabel metal3 s 31704 63388 31802 63486 4 gnd
port 3 nsew
rlabel metal3 s 29639 61839 29737 61937 4 vdd
port 2 nsew
rlabel metal3 s 30768 61248 30866 61346 4 vdd
port 2 nsew
rlabel metal3 s 32697 65911 32795 66009 4 vdd
port 2 nsew
rlabel metal3 s 32952 63388 33050 63486 4 gnd
port 3 nsew
rlabel metal3 s 29035 65137 29133 65235 4 gnd
port 3 nsew
rlabel metal3 s 27529 61839 27627 61937 4 vdd
port 2 nsew
rlabel metal3 s 27024 61248 27122 61346 4 vdd
port 2 nsew
rlabel metal3 s 31392 61248 31490 61346 4 vdd
port 2 nsew
rlabel metal3 s 26457 65911 26555 66009 4 vdd
port 2 nsew
rlabel metal3 s 32709 67071 32807 67169 4 gnd
port 3 nsew
rlabel metal3 s 27960 63388 28058 63486 4 gnd
port 3 nsew
rlabel metal3 s 30025 61839 30123 61937 4 vdd
port 2 nsew
rlabel metal3 s 25895 61839 25993 61937 4 vdd
port 2 nsew
rlabel metal3 s 30887 61839 30985 61937 4 vdd
port 2 nsew
rlabel metal3 s 27717 66749 27815 66847 4 vdd
port 2 nsew
rlabel metal3 s 26400 61248 26498 61346 4 vdd
port 2 nsew
rlabel metal3 s 25776 61248 25874 61346 4 vdd
port 2 nsew
rlabel metal3 s 28777 61839 28875 61937 4 vdd
port 2 nsew
rlabel metal3 s 31531 65137 31629 65235 4 gnd
port 3 nsew
rlabel metal3 s 28272 61248 28370 61346 4 vdd
port 2 nsew
rlabel metal3 s 29208 63388 29306 63486 4 gnd
port 3 nsew
rlabel metal3 s 27717 67071 27815 67169 4 gnd
port 3 nsew
rlabel metal3 s 26469 66749 26567 66847 4 vdd
port 2 nsew
rlabel metal3 s 26712 63388 26810 63486 4 gnd
port 3 nsew
rlabel metal3 s 31461 67071 31559 67169 4 gnd
port 3 nsew
rlabel metal3 s 31273 61839 31371 61937 4 vdd
port 2 nsew
rlabel metal3 s 26281 61839 26379 61937 4 vdd
port 2 nsew
rlabel metal3 s 27143 61839 27241 61937 4 vdd
port 2 nsew
rlabel metal3 s 26539 65137 26637 65235 4 gnd
port 3 nsew
rlabel metal3 s 30283 65137 30381 65235 4 gnd
port 3 nsew
rlabel metal3 s 28965 66749 29063 66847 4 vdd
port 2 nsew
rlabel metal3 s 28965 67071 29063 67169 4 gnd
port 3 nsew
rlabel metal3 s 30144 61248 30242 61346 4 vdd
port 2 nsew
rlabel metal3 s 27787 65137 27885 65235 4 gnd
port 3 nsew
rlabel metal3 s 30213 66749 30311 66847 4 vdd
port 2 nsew
rlabel metal3 s 33264 61248 33362 61346 4 vdd
port 2 nsew
rlabel metal3 s 33383 61839 33481 61937 4 vdd
port 2 nsew
rlabel metal3 s 30213 67071 30311 67169 4 gnd
port 3 nsew
rlabel metal3 s 31449 65911 31547 66009 4 vdd
port 2 nsew
rlabel metal3 s 28391 61839 28489 61937 4 vdd
port 2 nsew
rlabel metal3 s 32640 61248 32738 61346 4 vdd
port 2 nsew
rlabel metal3 s 32521 61839 32619 61937 4 vdd
port 2 nsew
rlabel metal3 s 30456 63388 30554 63486 4 gnd
port 3 nsew
rlabel metal3 s 31461 66749 31559 66847 4 vdd
port 2 nsew
rlabel metal3 s 27705 65911 27803 66009 4 vdd
port 2 nsew
rlabel metal3 s 27648 61248 27746 61346 4 vdd
port 2 nsew
rlabel metal3 s 26469 67071 26567 67169 4 gnd
port 3 nsew
rlabel metal3 s 32016 61248 32114 61346 4 vdd
port 2 nsew
rlabel metal3 s 28896 61248 28994 61346 4 vdd
port 2 nsew
rlabel metal3 s 29520 61248 29618 61346 4 vdd
port 2 nsew
rlabel metal3 s 30201 65911 30299 66009 4 vdd
port 2 nsew
rlabel metal3 s 32709 66749 32807 66847 4 vdd
port 2 nsew
rlabel metal3 s 25464 63388 25562 63486 4 gnd
port 3 nsew
rlabel metal3 s 22656 61248 22754 61346 4 vdd
port 2 nsew
rlabel metal3 s 25033 61839 25131 61937 4 vdd
port 2 nsew
rlabel metal3 s 17733 66749 17831 66847 4 vdd
port 2 nsew
rlabel metal3 s 17664 61248 17762 61346 4 vdd
port 2 nsew
rlabel metal3 s 25221 67071 25319 67169 4 gnd
port 3 nsew
rlabel metal3 s 23961 65911 24059 66009 4 vdd
port 2 nsew
rlabel metal3 s 18407 61839 18505 61937 4 vdd
port 2 nsew
rlabel metal3 s 23280 61248 23378 61346 4 vdd
port 2 nsew
rlabel metal3 s 21408 61248 21506 61346 4 vdd
port 2 nsew
rlabel metal3 s 19051 65137 19149 65235 4 gnd
port 3 nsew
rlabel metal3 s 19655 61839 19753 61937 4 vdd
port 2 nsew
rlabel metal3 s 20903 61839 21001 61937 4 vdd
port 2 nsew
rlabel metal3 s 20041 61839 20139 61937 4 vdd
port 2 nsew
rlabel metal3 s 21289 61839 21387 61937 4 vdd
port 2 nsew
rlabel metal3 s 18981 67071 19079 67169 4 gnd
port 3 nsew
rlabel metal3 s 17733 67071 17831 67169 4 gnd
port 3 nsew
rlabel metal3 s 25291 65137 25389 65235 4 gnd
port 3 nsew
rlabel metal3 s 17976 63388 18074 63486 4 gnd
port 3 nsew
rlabel metal3 s 23785 61839 23883 61937 4 vdd
port 2 nsew
rlabel metal3 s 18981 66749 19079 66847 4 vdd
port 2 nsew
rlabel metal3 s 18969 65911 19067 66009 4 vdd
port 2 nsew
rlabel metal3 s 25152 61248 25250 61346 4 vdd
port 2 nsew
rlabel metal3 s 24216 63388 24314 63486 4 gnd
port 3 nsew
rlabel metal3 s 21477 67071 21575 67169 4 gnd
port 3 nsew
rlabel metal3 s 18793 61839 18891 61937 4 vdd
port 2 nsew
rlabel metal3 s 21477 66749 21575 66847 4 vdd
port 2 nsew
rlabel metal3 s 20160 61248 20258 61346 4 vdd
port 2 nsew
rlabel metal3 s 20299 65137 20397 65235 4 gnd
port 3 nsew
rlabel metal3 s 24647 61839 24745 61937 4 vdd
port 2 nsew
rlabel metal3 s 19536 61248 19634 61346 4 vdd
port 2 nsew
rlabel metal3 s 23973 66749 24071 66847 4 vdd
port 2 nsew
rlabel metal3 s 21465 65911 21563 66009 4 vdd
port 2 nsew
rlabel metal3 s 22725 67071 22823 67169 4 gnd
port 3 nsew
rlabel metal3 s 21720 63388 21818 63486 4 gnd
port 3 nsew
rlabel metal3 s 23973 67071 24071 67169 4 gnd
port 3 nsew
rlabel metal3 s 25221 66749 25319 66847 4 vdd
port 2 nsew
rlabel metal3 s 22151 61839 22249 61937 4 vdd
port 2 nsew
rlabel metal3 s 18912 61248 19010 61346 4 vdd
port 2 nsew
rlabel metal3 s 19224 63388 19322 63486 4 gnd
port 3 nsew
rlabel metal3 s 22032 61248 22130 61346 4 vdd
port 2 nsew
rlabel metal3 s 18288 61248 18386 61346 4 vdd
port 2 nsew
rlabel metal3 s 22713 65911 22811 66009 4 vdd
port 2 nsew
rlabel metal3 s 23399 61839 23497 61937 4 vdd
port 2 nsew
rlabel metal3 s 23904 61248 24002 61346 4 vdd
port 2 nsew
rlabel metal3 s 22968 63388 23066 63486 4 gnd
port 3 nsew
rlabel metal3 s 21547 65137 21645 65235 4 gnd
port 3 nsew
rlabel metal3 s 22795 65137 22893 65235 4 gnd
port 3 nsew
rlabel metal3 s 17803 65137 17901 65235 4 gnd
port 3 nsew
rlabel metal3 s 24528 61248 24626 61346 4 vdd
port 2 nsew
rlabel metal3 s 20217 65911 20315 66009 4 vdd
port 2 nsew
rlabel metal3 s 24043 65137 24141 65235 4 gnd
port 3 nsew
rlabel metal3 s 25209 65911 25307 66009 4 vdd
port 2 nsew
rlabel metal3 s 22537 61839 22635 61937 4 vdd
port 2 nsew
rlabel metal3 s 22725 66749 22823 66847 4 vdd
port 2 nsew
rlabel metal3 s 20472 63388 20570 63486 4 gnd
port 3 nsew
rlabel metal3 s 17721 65911 17819 66009 4 vdd
port 2 nsew
rlabel metal3 s 20784 61248 20882 61346 4 vdd
port 2 nsew
rlabel metal3 s 17545 61839 17643 61937 4 vdd
port 2 nsew
rlabel metal3 s 20229 67071 20327 67169 4 gnd
port 3 nsew
rlabel metal3 s 20229 66749 20327 66847 4 vdd
port 2 nsew
rlabel metal3 s 13296 61248 13394 61346 4 vdd
port 2 nsew
rlabel metal3 s 13920 61248 14018 61346 4 vdd
port 2 nsew
rlabel metal3 s 13989 66749 14087 66847 4 vdd
port 2 nsew
rlabel metal3 s 15480 63388 15578 63486 4 gnd
port 3 nsew
rlabel metal3 s 12600 60134 12698 60232 4 gnd
port 3 nsew
rlabel metal3 s 12600 60687 12698 60785 4 gnd
port 3 nsew
rlabel metal3 s 16416 61248 16514 61346 4 vdd
port 2 nsew
rlabel metal3 s 16473 65911 16571 66009 4 vdd
port 2 nsew
rlabel metal3 s 15307 65137 15405 65235 4 gnd
port 3 nsew
rlabel metal3 s 16485 66749 16583 66847 4 vdd
port 2 nsew
rlabel metal3 s 14059 65137 14157 65235 4 gnd
port 3 nsew
rlabel metal3 s 12600 59344 12698 59442 4 gnd
port 3 nsew
rlabel metal3 s 14544 61248 14642 61346 4 vdd
port 2 nsew
rlabel metal3 s 17040 61248 17138 61346 4 vdd
port 2 nsew
rlabel metal3 s 13989 67071 14087 67169 4 gnd
port 3 nsew
rlabel metal3 s 15237 67071 15335 67169 4 gnd
port 3 nsew
rlabel metal3 s 12600 58870 12698 58968 4 gnd
port 3 nsew
rlabel metal3 s 13977 65911 14075 66009 4 vdd
port 2 nsew
rlabel metal3 s 12234 61034 12332 61132 4 gnd
port 3 nsew
rlabel metal3 s 12600 59660 12698 59758 4 gnd
port 3 nsew
rlabel metal3 s 12600 59897 12698 59995 4 gnd
port 3 nsew
rlabel metal3 s 15225 65911 15323 66009 4 vdd
port 2 nsew
rlabel metal3 s 12600 60450 12698 60548 4 gnd
port 3 nsew
rlabel metal3 s 14663 61839 14761 61937 4 vdd
port 2 nsew
rlabel metal3 s 15168 61248 15266 61346 4 vdd
port 2 nsew
rlabel metal3 s 16485 67071 16583 67169 4 gnd
port 3 nsew
rlabel metal3 s 16297 61839 16395 61937 4 vdd
port 2 nsew
rlabel metal3 s 15911 61839 16009 61937 4 vdd
port 2 nsew
rlabel metal3 s 15237 66749 15335 66847 4 vdd
port 2 nsew
rlabel metal3 s 12600 59107 12698 59205 4 gnd
port 3 nsew
rlabel metal3 s 16728 63388 16826 63486 4 gnd
port 3 nsew
rlabel metal3 s 16555 65137 16653 65235 4 gnd
port 3 nsew
rlabel metal3 s 13801 61839 13899 61937 4 vdd
port 2 nsew
rlabel metal3 s 17159 61839 17257 61937 4 vdd
port 2 nsew
rlabel metal3 s 14232 63388 14330 63486 4 gnd
port 3 nsew
rlabel metal3 s 15792 61248 15890 61346 4 vdd
port 2 nsew
rlabel metal3 s 15049 61839 15147 61937 4 vdd
port 2 nsew
rlabel metal3 s 7264 59502 7362 59600 4 gnd
port 3 nsew
rlabel metal3 s 6025 60315 6123 60413 4 gnd
port 3 nsew
rlabel metal3 s 6882 59883 6980 59981 4 vdd
port 2 nsew
rlabel metal3 s 6025 59525 6123 59623 4 gnd
port 3 nsew
rlabel metal3 s 7264 58712 7362 58810 4 gnd
port 3 nsew
rlabel metal3 s 7264 60292 7362 60390 4 gnd
port 3 nsew
rlabel metal3 s 6450 60315 6548 60413 4 vdd
port 2 nsew
rlabel metal3 s 6450 59093 6548 59191 4 vdd
port 2 nsew
rlabel metal3 s 6882 59525 6980 59623 4 vdd
port 2 nsew
rlabel metal3 s 6882 60315 6980 60413 4 vdd
port 2 nsew
rlabel metal3 s 6025 59941 6123 60039 4 gnd
port 3 nsew
rlabel metal3 s 6882 59093 6980 59191 4 vdd
port 2 nsew
rlabel metal3 s 6025 59151 6123 59249 4 gnd
port 3 nsew
rlabel metal3 s 7264 59107 7362 59205 4 gnd
port 3 nsew
rlabel metal3 s 7660 59107 7758 59205 4 vdd
port 2 nsew
rlabel metal3 s 6025 58735 6123 58833 4 gnd
port 3 nsew
rlabel metal3 s 6450 59525 6548 59623 4 vdd
port 2 nsew
rlabel metal3 s 7660 59502 7758 59600 4 vdd
port 2 nsew
rlabel metal3 s 7660 60292 7758 60390 4 vdd
port 2 nsew
rlabel metal3 s 6882 58735 6980 58833 4 vdd
port 2 nsew
rlabel metal3 s 7264 59897 7362 59995 4 gnd
port 3 nsew
rlabel metal3 s 6450 58735 6548 58833 4 vdd
port 2 nsew
rlabel metal3 s 7660 58712 7758 58810 4 vdd
port 2 nsew
rlabel metal3 s 6450 59883 6548 59981 4 vdd
port 2 nsew
rlabel metal3 s 7660 59897 7758 59995 4 vdd
port 2 nsew
rlabel metal3 s 7264 55947 7362 56045 4 gnd
port 3 nsew
rlabel metal3 s 7264 56737 7362 56835 4 gnd
port 3 nsew
rlabel metal3 s 6882 57513 6980 57611 4 vdd
port 2 nsew
rlabel metal3 s 6025 58361 6123 58459 4 gnd
port 3 nsew
rlabel metal3 s 7660 56737 7758 56835 4 vdd
port 2 nsew
rlabel metal3 s 6450 54785 6548 54883 4 vdd
port 2 nsew
rlabel metal3 s 6450 57945 6548 58043 4 vdd
port 2 nsew
rlabel metal3 s 6025 56781 6123 56879 4 gnd
port 3 nsew
rlabel metal3 s 6025 55991 6123 56089 4 gnd
port 3 nsew
rlabel metal3 s 6882 56365 6980 56463 4 vdd
port 2 nsew
rlabel metal3 s 6450 57513 6548 57611 4 vdd
port 2 nsew
rlabel metal3 s 7264 54762 7362 54860 4 gnd
port 3 nsew
rlabel metal3 s 6025 55201 6123 55299 4 gnd
port 3 nsew
rlabel metal3 s 6450 57155 6548 57253 4 vdd
port 2 nsew
rlabel metal3 s 7660 56342 7758 56440 4 vdd
port 2 nsew
rlabel metal3 s 6450 56365 6548 56463 4 vdd
port 2 nsew
rlabel metal3 s 6450 55575 6548 55673 4 vdd
port 2 nsew
rlabel metal3 s 6025 56365 6123 56463 4 gnd
port 3 nsew
rlabel metal3 s 7660 57132 7758 57230 4 vdd
port 2 nsew
rlabel metal3 s 7660 57527 7758 57625 4 vdd
port 2 nsew
rlabel metal3 s 7264 57922 7362 58020 4 gnd
port 3 nsew
rlabel metal3 s 6450 55143 6548 55241 4 vdd
port 2 nsew
rlabel metal3 s 7264 57132 7362 57230 4 gnd
port 3 nsew
rlabel metal3 s 6025 57945 6123 58043 4 gnd
port 3 nsew
rlabel metal3 s 6882 55933 6980 56031 4 vdd
port 2 nsew
rlabel metal3 s 6450 55933 6548 56031 4 vdd
port 2 nsew
rlabel metal3 s 6882 57945 6980 58043 4 vdd
port 2 nsew
rlabel metal3 s 7264 58317 7362 58415 4 gnd
port 3 nsew
rlabel metal3 s 6882 57155 6980 57253 4 vdd
port 2 nsew
rlabel metal3 s 7660 55157 7758 55255 4 vdd
port 2 nsew
rlabel metal3 s 7264 56342 7362 56440 4 gnd
port 3 nsew
rlabel metal3 s 7264 57527 7362 57625 4 gnd
port 3 nsew
rlabel metal3 s 6025 57155 6123 57253 4 gnd
port 3 nsew
rlabel metal3 s 6025 54785 6123 54883 4 gnd
port 3 nsew
rlabel metal3 s 6025 55575 6123 55673 4 gnd
port 3 nsew
rlabel metal3 s 6882 55143 6980 55241 4 vdd
port 2 nsew
rlabel metal3 s 6882 56723 6980 56821 4 vdd
port 2 nsew
rlabel metal3 s 6882 55575 6980 55673 4 vdd
port 2 nsew
rlabel metal3 s 7660 55552 7758 55650 4 vdd
port 2 nsew
rlabel metal3 s 7660 57922 7758 58020 4 vdd
port 2 nsew
rlabel metal3 s 7660 58317 7758 58415 4 vdd
port 2 nsew
rlabel metal3 s 6882 54785 6980 54883 4 vdd
port 2 nsew
rlabel metal3 s 7660 54762 7758 54860 4 vdd
port 2 nsew
rlabel metal3 s 6450 56723 6548 56821 4 vdd
port 2 nsew
rlabel metal3 s 6450 58303 6548 58401 4 vdd
port 2 nsew
rlabel metal3 s 7264 55157 7362 55255 4 gnd
port 3 nsew
rlabel metal3 s 7264 55552 7362 55650 4 gnd
port 3 nsew
rlabel metal3 s 6882 58303 6980 58401 4 vdd
port 2 nsew
rlabel metal3 s 6025 57571 6123 57669 4 gnd
port 3 nsew
rlabel metal3 s 7660 55947 7758 56045 4 vdd
port 2 nsew
rlabel metal3 s 7264 51997 7362 52095 4 gnd
port 3 nsew
rlabel metal3 s 6450 51983 6548 52081 4 vdd
port 2 nsew
rlabel metal3 s 6882 52773 6980 52871 4 vdd
port 2 nsew
rlabel metal3 s 6882 51193 6980 51291 4 vdd
port 2 nsew
rlabel metal3 s 6450 53995 6548 54093 4 vdd
port 2 nsew
rlabel metal3 s 7660 52787 7758 52885 4 vdd
port 2 nsew
rlabel metal3 s 6025 51251 6123 51349 4 gnd
port 3 nsew
rlabel metal3 s 6882 50403 6980 50501 4 vdd
port 2 nsew
rlabel metal3 s 7264 50417 7362 50515 4 gnd
port 3 nsew
rlabel metal3 s 6882 50835 6980 50933 4 vdd
port 2 nsew
rlabel metal3 s 6882 51625 6980 51723 4 vdd
port 2 nsew
rlabel metal3 s 6450 51193 6548 51291 4 vdd
port 2 nsew
rlabel metal3 s 7264 51207 7362 51305 4 gnd
port 3 nsew
rlabel metal3 s 7660 53972 7758 54070 4 vdd
port 2 nsew
rlabel metal3 s 6025 54411 6123 54509 4 gnd
port 3 nsew
rlabel metal3 s 6025 50461 6123 50559 4 gnd
port 3 nsew
rlabel metal3 s 6882 53563 6980 53661 4 vdd
port 2 nsew
rlabel metal3 s 7660 53182 7758 53280 4 vdd
port 2 nsew
rlabel metal3 s 6450 50835 6548 50933 4 vdd
port 2 nsew
rlabel metal3 s 6882 51983 6980 52081 4 vdd
port 2 nsew
rlabel metal3 s 7660 52392 7758 52490 4 vdd
port 2 nsew
rlabel metal3 s 7264 53972 7362 54070 4 gnd
port 3 nsew
rlabel metal3 s 6882 52415 6980 52513 4 vdd
port 2 nsew
rlabel metal3 s 7660 51997 7758 52095 4 vdd
port 2 nsew
rlabel metal3 s 6025 52041 6123 52139 4 gnd
port 3 nsew
rlabel metal3 s 6882 54353 6980 54451 4 vdd
port 2 nsew
rlabel metal3 s 6025 52831 6123 52929 4 gnd
port 3 nsew
rlabel metal3 s 6450 53563 6548 53661 4 vdd
port 2 nsew
rlabel metal3 s 7660 51207 7758 51305 4 vdd
port 2 nsew
rlabel metal3 s 7264 52787 7362 52885 4 gnd
port 3 nsew
rlabel metal3 s 6025 53205 6123 53303 4 gnd
port 3 nsew
rlabel metal3 s 6882 53205 6980 53303 4 vdd
port 2 nsew
rlabel metal3 s 7660 54367 7758 54465 4 vdd
port 2 nsew
rlabel metal3 s 6025 52415 6123 52513 4 gnd
port 3 nsew
rlabel metal3 s 6025 53995 6123 54093 4 gnd
port 3 nsew
rlabel metal3 s 7660 50812 7758 50910 4 vdd
port 2 nsew
rlabel metal3 s 6450 52415 6548 52513 4 vdd
port 2 nsew
rlabel metal3 s 7264 52392 7362 52490 4 gnd
port 3 nsew
rlabel metal3 s 6882 53995 6980 54093 4 vdd
port 2 nsew
rlabel metal3 s 7264 53182 7362 53280 4 gnd
port 3 nsew
rlabel metal3 s 6450 53205 6548 53303 4 vdd
port 2 nsew
rlabel metal3 s 7264 50812 7362 50910 4 gnd
port 3 nsew
rlabel metal3 s 7660 51602 7758 51700 4 vdd
port 2 nsew
rlabel metal3 s 6450 54353 6548 54451 4 vdd
port 2 nsew
rlabel metal3 s 7660 53577 7758 53675 4 vdd
port 2 nsew
rlabel metal3 s 7660 50417 7758 50515 4 vdd
port 2 nsew
rlabel metal3 s 6025 53621 6123 53719 4 gnd
port 3 nsew
rlabel metal3 s 6450 50403 6548 50501 4 vdd
port 2 nsew
rlabel metal3 s 7264 51602 7362 51700 4 gnd
port 3 nsew
rlabel metal3 s 7264 54367 7362 54465 4 gnd
port 3 nsew
rlabel metal3 s 7264 53577 7362 53675 4 gnd
port 3 nsew
rlabel metal3 s 6450 51625 6548 51723 4 vdd
port 2 nsew
rlabel metal3 s 6025 51625 6123 51723 4 gnd
port 3 nsew
rlabel metal3 s 6450 52773 6548 52871 4 vdd
port 2 nsew
rlabel metal3 s 6025 50835 6123 50933 4 gnd
port 3 nsew
rlabel metal3 s 12600 57527 12698 57625 4 gnd
port 3 nsew
rlabel metal3 s 12600 52550 12698 52648 4 gnd
port 3 nsew
rlabel metal3 s 12600 51444 12698 51542 4 gnd
port 3 nsew
rlabel metal3 s 12600 55157 12698 55255 4 gnd
port 3 nsew
rlabel metal3 s 12600 53577 12698 53675 4 gnd
port 3 nsew
rlabel metal3 s 12600 55394 12698 55492 4 gnd
port 3 nsew
rlabel metal3 s 12600 57290 12698 57388 4 gnd
port 3 nsew
rlabel metal3 s 12600 56737 12698 56835 4 gnd
port 3 nsew
rlabel metal3 s 12600 51997 12698 52095 4 gnd
port 3 nsew
rlabel metal3 s 12600 52234 12698 52332 4 gnd
port 3 nsew
rlabel metal3 s 12600 50970 12698 51068 4 gnd
port 3 nsew
rlabel metal3 s 12600 54920 12698 55018 4 gnd
port 3 nsew
rlabel metal3 s 12600 58554 12698 58652 4 gnd
port 3 nsew
rlabel metal3 s 12600 51760 12698 51858 4 gnd
port 3 nsew
rlabel metal3 s 12600 54604 12698 54702 4 gnd
port 3 nsew
rlabel metal3 s 12600 52787 12698 52885 4 gnd
port 3 nsew
rlabel metal3 s 12600 53814 12698 53912 4 gnd
port 3 nsew
rlabel metal3 s 12600 57764 12698 57862 4 gnd
port 3 nsew
rlabel metal3 s 12600 55947 12698 56045 4 gnd
port 3 nsew
rlabel metal3 s 12600 54367 12698 54465 4 gnd
port 3 nsew
rlabel metal3 s 12600 51207 12698 51305 4 gnd
port 3 nsew
rlabel metal3 s 12600 58317 12698 58415 4 gnd
port 3 nsew
rlabel metal3 s 12600 53024 12698 53122 4 gnd
port 3 nsew
rlabel metal3 s 12600 53340 12698 53438 4 gnd
port 3 nsew
rlabel metal3 s 12600 58080 12698 58178 4 gnd
port 3 nsew
rlabel metal3 s 12600 56974 12698 57072 4 gnd
port 3 nsew
rlabel metal3 s 12600 54130 12698 54228 4 gnd
port 3 nsew
rlabel metal3 s 12600 56500 12698 56598 4 gnd
port 3 nsew
rlabel metal3 s 12600 50654 12698 50752 4 gnd
port 3 nsew
rlabel metal3 s 12600 50417 12698 50515 4 gnd
port 3 nsew
rlabel metal3 s 12600 55710 12698 55808 4 gnd
port 3 nsew
rlabel metal3 s 12600 56184 12698 56282 4 gnd
port 3 nsew
rlabel metal3 s 12600 43544 12698 43642 4 gnd
port 3 nsew
rlabel metal3 s 12600 42280 12698 42378 4 gnd
port 3 nsew
rlabel metal3 s 12600 47020 12698 47118 4 gnd
port 3 nsew
rlabel metal3 s 12600 43070 12698 43168 4 gnd
port 3 nsew
rlabel metal3 s 12600 41964 12698 42062 4 gnd
port 3 nsew
rlabel metal3 s 12600 49627 12698 49725 4 gnd
port 3 nsew
rlabel metal3 s 12600 43860 12698 43958 4 gnd
port 3 nsew
rlabel metal3 s 12600 44097 12698 44195 4 gnd
port 3 nsew
rlabel metal3 s 12600 42754 12698 42852 4 gnd
port 3 nsew
rlabel metal3 s 12600 44887 12698 44985 4 gnd
port 3 nsew
rlabel metal3 s 12600 47494 12698 47592 4 gnd
port 3 nsew
rlabel metal3 s 12600 45440 12698 45538 4 gnd
port 3 nsew
rlabel metal3 s 12600 49864 12698 49962 4 gnd
port 3 nsew
rlabel metal3 s 12600 50180 12698 50278 4 gnd
port 3 nsew
rlabel metal3 s 12600 48600 12698 48698 4 gnd
port 3 nsew
rlabel metal3 s 12600 45914 12698 46012 4 gnd
port 3 nsew
rlabel metal3 s 12600 46704 12698 46802 4 gnd
port 3 nsew
rlabel metal3 s 12600 42517 12698 42615 4 gnd
port 3 nsew
rlabel metal3 s 12600 48284 12698 48382 4 gnd
port 3 nsew
rlabel metal3 s 12600 48047 12698 48145 4 gnd
port 3 nsew
rlabel metal3 s 12600 49390 12698 49488 4 gnd
port 3 nsew
rlabel metal3 s 12600 47810 12698 47908 4 gnd
port 3 nsew
rlabel metal3 s 12600 49074 12698 49172 4 gnd
port 3 nsew
rlabel metal3 s 12600 47257 12698 47355 4 gnd
port 3 nsew
rlabel metal3 s 12600 46230 12698 46328 4 gnd
port 3 nsew
rlabel metal3 s 12600 45124 12698 45222 4 gnd
port 3 nsew
rlabel metal3 s 12600 45677 12698 45775 4 gnd
port 3 nsew
rlabel metal3 s 12600 48837 12698 48935 4 gnd
port 3 nsew
rlabel metal3 s 12600 44650 12698 44748 4 gnd
port 3 nsew
rlabel metal3 s 12600 43307 12698 43405 4 gnd
port 3 nsew
rlabel metal3 s 12600 46467 12698 46565 4 gnd
port 3 nsew
rlabel metal3 s 12600 44334 12698 44432 4 gnd
port 3 nsew
rlabel metal3 s 6450 46453 6548 46551 4 vdd
port 2 nsew
rlabel metal3 s 6882 49613 6980 49711 4 vdd
port 2 nsew
rlabel metal3 s 6450 48033 6548 48131 4 vdd
port 2 nsew
rlabel metal3 s 7660 49627 7758 49725 4 vdd
port 2 nsew
rlabel metal3 s 6450 47243 6548 47341 4 vdd
port 2 nsew
rlabel metal3 s 7660 50022 7758 50120 4 vdd
port 2 nsew
rlabel metal3 s 6025 48091 6123 48189 4 gnd
port 3 nsew
rlabel metal3 s 6882 46453 6980 46551 4 vdd
port 2 nsew
rlabel metal3 s 6025 50045 6123 50143 4 gnd
port 3 nsew
rlabel metal3 s 6882 47243 6980 47341 4 vdd
port 2 nsew
rlabel metal3 s 7660 47257 7758 47355 4 vdd
port 2 nsew
rlabel metal3 s 6450 48823 6548 48921 4 vdd
port 2 nsew
rlabel metal3 s 6450 48465 6548 48563 4 vdd
port 2 nsew
rlabel metal3 s 6882 48823 6980 48921 4 vdd
port 2 nsew
rlabel metal3 s 6882 48465 6980 48563 4 vdd
port 2 nsew
rlabel metal3 s 7264 48047 7362 48145 4 gnd
port 3 nsew
rlabel metal3 s 6025 46511 6123 46609 4 gnd
port 3 nsew
rlabel metal3 s 6882 48033 6980 48131 4 vdd
port 2 nsew
rlabel metal3 s 7264 49627 7362 49725 4 gnd
port 3 nsew
rlabel metal3 s 6025 48881 6123 48979 4 gnd
port 3 nsew
rlabel metal3 s 6882 47675 6980 47773 4 vdd
port 2 nsew
rlabel metal3 s 7660 47652 7758 47750 4 vdd
port 2 nsew
rlabel metal3 s 7264 48442 7362 48540 4 gnd
port 3 nsew
rlabel metal3 s 6450 49613 6548 49711 4 vdd
port 2 nsew
rlabel metal3 s 7264 47257 7362 47355 4 gnd
port 3 nsew
rlabel metal3 s 6882 46885 6980 46983 4 vdd
port 2 nsew
rlabel metal3 s 7264 48837 7362 48935 4 gnd
port 3 nsew
rlabel metal3 s 6450 50045 6548 50143 4 vdd
port 2 nsew
rlabel metal3 s 7660 46862 7758 46960 4 vdd
port 2 nsew
rlabel metal3 s 7264 47652 7362 47750 4 gnd
port 3 nsew
rlabel metal3 s 7264 46862 7362 46960 4 gnd
port 3 nsew
rlabel metal3 s 6025 49671 6123 49769 4 gnd
port 3 nsew
rlabel metal3 s 7264 50022 7362 50120 4 gnd
port 3 nsew
rlabel metal3 s 7264 49232 7362 49330 4 gnd
port 3 nsew
rlabel metal3 s 6882 50045 6980 50143 4 vdd
port 2 nsew
rlabel metal3 s 7660 48442 7758 48540 4 vdd
port 2 nsew
rlabel metal3 s 6882 49255 6980 49353 4 vdd
port 2 nsew
rlabel metal3 s 6025 47301 6123 47399 4 gnd
port 3 nsew
rlabel metal3 s 7660 49232 7758 49330 4 vdd
port 2 nsew
rlabel metal3 s 6025 48465 6123 48563 4 gnd
port 3 nsew
rlabel metal3 s 7264 46467 7362 46565 4 gnd
port 3 nsew
rlabel metal3 s 7660 48047 7758 48145 4 vdd
port 2 nsew
rlabel metal3 s 6025 49255 6123 49353 4 gnd
port 3 nsew
rlabel metal3 s 6025 47675 6123 47773 4 gnd
port 3 nsew
rlabel metal3 s 7660 46467 7758 46565 4 vdd
port 2 nsew
rlabel metal3 s 6450 46885 6548 46983 4 vdd
port 2 nsew
rlabel metal3 s 6450 47675 6548 47773 4 vdd
port 2 nsew
rlabel metal3 s 6450 49255 6548 49353 4 vdd
port 2 nsew
rlabel metal3 s 6025 46885 6123 46983 4 gnd
port 3 nsew
rlabel metal3 s 7660 48837 7758 48935 4 vdd
port 2 nsew
rlabel metal3 s 7660 44887 7758 44985 4 vdd
port 2 nsew
rlabel metal3 s 6882 46095 6980 46193 4 vdd
port 2 nsew
rlabel metal3 s 7264 43702 7362 43800 4 gnd
port 3 nsew
rlabel metal3 s 6450 44873 6548 44971 4 vdd
port 2 nsew
rlabel metal3 s 7264 42517 7362 42615 4 gnd
port 3 nsew
rlabel metal3 s 7660 43307 7758 43405 4 vdd
port 2 nsew
rlabel metal3 s 7660 42122 7758 42220 4 vdd
port 2 nsew
rlabel metal3 s 7660 45677 7758 45775 4 vdd
port 2 nsew
rlabel metal3 s 6025 44931 6123 45029 4 gnd
port 3 nsew
rlabel metal3 s 6450 45305 6548 45403 4 vdd
port 2 nsew
rlabel metal3 s 6882 44873 6980 44971 4 vdd
port 2 nsew
rlabel metal3 s 7264 44097 7362 44195 4 gnd
port 3 nsew
rlabel metal3 s 7264 45677 7362 45775 4 gnd
port 3 nsew
rlabel metal3 s 6882 42503 6980 42601 4 vdd
port 2 nsew
rlabel metal3 s 6450 46095 6548 46193 4 vdd
port 2 nsew
rlabel metal3 s 7264 43307 7362 43405 4 gnd
port 3 nsew
rlabel metal3 s 6025 42145 6123 42243 4 gnd
port 3 nsew
rlabel metal3 s 6450 42503 6548 42601 4 vdd
port 2 nsew
rlabel metal3 s 6882 42935 6980 43033 4 vdd
port 2 nsew
rlabel metal3 s 6882 44515 6980 44613 4 vdd
port 2 nsew
rlabel metal3 s 7264 46072 7362 46170 4 gnd
port 3 nsew
rlabel metal3 s 7264 45282 7362 45380 4 gnd
port 3 nsew
rlabel metal3 s 7660 44492 7758 44590 4 vdd
port 2 nsew
rlabel metal3 s 7264 44492 7362 44590 4 gnd
port 3 nsew
rlabel metal3 s 6450 43725 6548 43823 4 vdd
port 2 nsew
rlabel metal3 s 6025 45305 6123 45403 4 gnd
port 3 nsew
rlabel metal3 s 6025 44515 6123 44613 4 gnd
port 3 nsew
rlabel metal3 s 6025 44141 6123 44239 4 gnd
port 3 nsew
rlabel metal3 s 6025 45721 6123 45819 4 gnd
port 3 nsew
rlabel metal3 s 7264 44887 7362 44985 4 gnd
port 3 nsew
rlabel metal3 s 6882 45663 6980 45761 4 vdd
port 2 nsew
rlabel metal3 s 6450 42145 6548 42243 4 vdd
port 2 nsew
rlabel metal3 s 6025 42935 6123 43033 4 gnd
port 3 nsew
rlabel metal3 s 6450 42935 6548 43033 4 vdd
port 2 nsew
rlabel metal3 s 6450 45663 6548 45761 4 vdd
port 2 nsew
rlabel metal3 s 6882 43293 6980 43391 4 vdd
port 2 nsew
rlabel metal3 s 6882 44083 6980 44181 4 vdd
port 2 nsew
rlabel metal3 s 6025 42561 6123 42659 4 gnd
port 3 nsew
rlabel metal3 s 7660 43702 7758 43800 4 vdd
port 2 nsew
rlabel metal3 s 6450 44083 6548 44181 4 vdd
port 2 nsew
rlabel metal3 s 7264 42122 7362 42220 4 gnd
port 3 nsew
rlabel metal3 s 6882 43725 6980 43823 4 vdd
port 2 nsew
rlabel metal3 s 6882 45305 6980 45403 4 vdd
port 2 nsew
rlabel metal3 s 6025 43351 6123 43449 4 gnd
port 3 nsew
rlabel metal3 s 6025 43725 6123 43823 4 gnd
port 3 nsew
rlabel metal3 s 7660 44097 7758 44195 4 vdd
port 2 nsew
rlabel metal3 s 7660 42912 7758 43010 4 vdd
port 2 nsew
rlabel metal3 s 6450 43293 6548 43391 4 vdd
port 2 nsew
rlabel metal3 s 7660 42517 7758 42615 4 vdd
port 2 nsew
rlabel metal3 s 7660 46072 7758 46170 4 vdd
port 2 nsew
rlabel metal3 s 7660 45282 7758 45380 4 vdd
port 2 nsew
rlabel metal3 s 6450 44515 6548 44613 4 vdd
port 2 nsew
rlabel metal3 s 6882 42145 6980 42243 4 vdd
port 2 nsew
rlabel metal3 s 7264 42912 7362 43010 4 gnd
port 3 nsew
rlabel metal3 s 6025 46095 6123 46193 4 gnd
port 3 nsew
rlabel metal3 s 6882 38985 6980 39083 4 vdd
port 2 nsew
rlabel metal3 s 6882 38553 6980 38651 4 vdd
port 2 nsew
rlabel metal3 s 6882 41355 6980 41453 4 vdd
port 2 nsew
rlabel metal3 s 6025 38985 6123 39083 4 gnd
port 3 nsew
rlabel metal3 s 7660 38962 7758 39060 4 vdd
port 2 nsew
rlabel metal3 s 6025 39775 6123 39873 4 gnd
port 3 nsew
rlabel metal3 s 7660 41727 7758 41825 4 vdd
port 2 nsew
rlabel metal3 s 6025 41771 6123 41869 4 gnd
port 3 nsew
rlabel metal3 s 7660 37777 7758 37875 4 vdd
port 2 nsew
rlabel metal3 s 7264 38962 7362 39060 4 gnd
port 3 nsew
rlabel metal3 s 7264 40542 7362 40640 4 gnd
port 3 nsew
rlabel metal3 s 6882 40565 6980 40663 4 vdd
port 2 nsew
rlabel metal3 s 7660 38567 7758 38665 4 vdd
port 2 nsew
rlabel metal3 s 6025 40191 6123 40289 4 gnd
port 3 nsew
rlabel metal3 s 6882 39775 6980 39873 4 vdd
port 2 nsew
rlabel metal3 s 6450 40133 6548 40231 4 vdd
port 2 nsew
rlabel metal3 s 7660 40937 7758 41035 4 vdd
port 2 nsew
rlabel metal3 s 6882 41713 6980 41811 4 vdd
port 2 nsew
rlabel metal3 s 7264 40147 7362 40245 4 gnd
port 3 nsew
rlabel metal3 s 6882 38195 6980 38293 4 vdd
port 2 nsew
rlabel metal3 s 6450 40923 6548 41021 4 vdd
port 2 nsew
rlabel metal3 s 6450 37763 6548 37861 4 vdd
port 2 nsew
rlabel metal3 s 6025 40565 6123 40663 4 gnd
port 3 nsew
rlabel metal3 s 7264 41332 7362 41430 4 gnd
port 3 nsew
rlabel metal3 s 7264 38172 7362 38270 4 gnd
port 3 nsew
rlabel metal3 s 6450 41713 6548 41811 4 vdd
port 2 nsew
rlabel metal3 s 6450 40565 6548 40663 4 vdd
port 2 nsew
rlabel metal3 s 7660 40542 7758 40640 4 vdd
port 2 nsew
rlabel metal3 s 6882 39343 6980 39441 4 vdd
port 2 nsew
rlabel metal3 s 6025 38195 6123 38293 4 gnd
port 3 nsew
rlabel metal3 s 6025 38611 6123 38709 4 gnd
port 3 nsew
rlabel metal3 s 6882 37763 6980 37861 4 vdd
port 2 nsew
rlabel metal3 s 7660 38172 7758 38270 4 vdd
port 2 nsew
rlabel metal3 s 6450 38985 6548 39083 4 vdd
port 2 nsew
rlabel metal3 s 6450 39343 6548 39441 4 vdd
port 2 nsew
rlabel metal3 s 6450 41355 6548 41453 4 vdd
port 2 nsew
rlabel metal3 s 6450 38195 6548 38293 4 vdd
port 2 nsew
rlabel metal3 s 6450 39775 6548 39873 4 vdd
port 2 nsew
rlabel metal3 s 7264 39752 7362 39850 4 gnd
port 3 nsew
rlabel metal3 s 7660 39357 7758 39455 4 vdd
port 2 nsew
rlabel metal3 s 7264 40937 7362 41035 4 gnd
port 3 nsew
rlabel metal3 s 7660 41332 7758 41430 4 vdd
port 2 nsew
rlabel metal3 s 6882 40923 6980 41021 4 vdd
port 2 nsew
rlabel metal3 s 6882 40133 6980 40231 4 vdd
port 2 nsew
rlabel metal3 s 7264 37777 7362 37875 4 gnd
port 3 nsew
rlabel metal3 s 7264 39357 7362 39455 4 gnd
port 3 nsew
rlabel metal3 s 6025 41355 6123 41453 4 gnd
port 3 nsew
rlabel metal3 s 7660 40147 7758 40245 4 vdd
port 2 nsew
rlabel metal3 s 6025 37821 6123 37919 4 gnd
port 3 nsew
rlabel metal3 s 6025 39401 6123 39499 4 gnd
port 3 nsew
rlabel metal3 s 7660 39752 7758 39850 4 vdd
port 2 nsew
rlabel metal3 s 7264 41727 7362 41825 4 gnd
port 3 nsew
rlabel metal3 s 7264 38567 7362 38665 4 gnd
port 3 nsew
rlabel metal3 s 6025 40981 6123 41079 4 gnd
port 3 nsew
rlabel metal3 s 6450 38553 6548 38651 4 vdd
port 2 nsew
rlabel metal3 s 7264 34617 7362 34715 4 gnd
port 3 nsew
rlabel metal3 s 8517 35391 8615 35489 4 vdd
port 2 nsew
rlabel metal3 s 7660 36197 7758 36295 4 vdd
port 2 nsew
rlabel metal3 s 6025 35825 6123 35923 4 gnd
port 3 nsew
rlabel metal3 s 7660 37382 7758 37480 4 vdd
port 2 nsew
rlabel metal3 s 6450 36183 6548 36281 4 vdd
port 2 nsew
rlabel metal3 s 6882 34603 6980 34701 4 vdd
port 2 nsew
rlabel metal3 s 7660 34617 7758 34715 4 vdd
port 2 nsew
rlabel metal3 s 6882 35825 6980 35923 4 vdd
port 2 nsew
rlabel metal3 s 6025 36615 6123 36713 4 gnd
port 3 nsew
rlabel metal3 s 7660 35407 7758 35505 4 vdd
port 2 nsew
rlabel metal3 s 6450 35393 6548 35491 4 vdd
port 2 nsew
rlabel metal3 s 7264 33827 7362 33925 4 gnd
port 3 nsew
rlabel metal3 s 7264 37382 7362 37480 4 gnd
port 3 nsew
rlabel metal3 s 7660 35012 7758 35110 4 vdd
port 2 nsew
rlabel metal3 s 6025 35035 6123 35133 4 gnd
port 3 nsew
rlabel metal3 s 7660 34222 7758 34320 4 vdd
port 2 nsew
rlabel metal3 s 6882 36973 6980 37071 4 vdd
port 2 nsew
rlabel metal3 s 6025 34245 6123 34343 4 gnd
port 3 nsew
rlabel metal3 s 6025 34661 6123 34759 4 gnd
port 3 nsew
rlabel metal3 s 6025 35451 6123 35549 4 gnd
port 3 nsew
rlabel metal3 s 6882 33813 6980 33911 4 vdd
port 2 nsew
rlabel metal3 s 7264 36197 7362 36295 4 gnd
port 3 nsew
rlabel metal3 s 6882 36183 6980 36281 4 vdd
port 2 nsew
rlabel metal3 s 6882 37405 6980 37503 4 vdd
port 2 nsew
rlabel metal3 s 6025 37031 6123 37129 4 gnd
port 3 nsew
rlabel metal3 s 6882 35035 6980 35133 4 vdd
port 2 nsew
rlabel metal3 s 7264 36987 7362 37085 4 gnd
port 3 nsew
rlabel metal3 s 6025 37405 6123 37503 4 gnd
port 3 nsew
rlabel metal3 s 6450 36973 6548 37071 4 vdd
port 2 nsew
rlabel metal3 s 7660 36987 7758 37085 4 vdd
port 2 nsew
rlabel metal3 s 6450 36615 6548 36713 4 vdd
port 2 nsew
rlabel metal3 s 7264 34222 7362 34320 4 gnd
port 3 nsew
rlabel metal3 s 6882 34245 6980 34343 4 vdd
port 2 nsew
rlabel metal3 s 6882 35393 6980 35491 4 vdd
port 2 nsew
rlabel metal3 s 7660 35802 7758 35900 4 vdd
port 2 nsew
rlabel metal3 s 6450 34603 6548 34701 4 vdd
port 2 nsew
rlabel metal3 s 6025 36241 6123 36339 4 gnd
port 3 nsew
rlabel metal3 s 6450 37405 6548 37503 4 vdd
port 2 nsew
rlabel metal3 s 6450 33813 6548 33911 4 vdd
port 2 nsew
rlabel metal3 s 7660 33827 7758 33925 4 vdd
port 2 nsew
rlabel metal3 s 8092 35392 8190 35490 4 gnd
port 3 nsew
rlabel metal3 s 7660 36592 7758 36690 4 vdd
port 2 nsew
rlabel metal3 s 6025 33871 6123 33969 4 gnd
port 3 nsew
rlabel metal3 s 7264 35802 7362 35900 4 gnd
port 3 nsew
rlabel metal3 s 6450 35825 6548 35923 4 vdd
port 2 nsew
rlabel metal3 s 7264 35012 7362 35110 4 gnd
port 3 nsew
rlabel metal3 s 6882 36615 6980 36713 4 vdd
port 2 nsew
rlabel metal3 s 6450 35035 6548 35133 4 vdd
port 2 nsew
rlabel metal3 s 7264 35407 7362 35505 4 gnd
port 3 nsew
rlabel metal3 s 6450 34245 6548 34343 4 vdd
port 2 nsew
rlabel metal3 s 7264 36592 7362 36690 4 gnd
port 3 nsew
rlabel metal3 s 12600 40937 12698 41035 4 gnd
port 3 nsew
rlabel metal3 s 12600 41490 12698 41588 4 gnd
port 3 nsew
rlabel metal3 s 12600 33590 12698 33688 4 gnd
port 3 nsew
rlabel metal3 s 12600 36750 12698 36848 4 gnd
port 3 nsew
rlabel metal3 s 12600 37224 12698 37322 4 gnd
port 3 nsew
rlabel metal3 s 12600 39357 12698 39455 4 gnd
port 3 nsew
rlabel metal3 s 12600 38567 12698 38665 4 gnd
port 3 nsew
rlabel metal3 s 12600 33827 12698 33925 4 gnd
port 3 nsew
rlabel metal3 s 12600 38014 12698 38112 4 gnd
port 3 nsew
rlabel metal3 s 12600 39594 12698 39692 4 gnd
port 3 nsew
rlabel metal3 s 11208 35407 11306 35505 4 vdd
port 2 nsew
rlabel metal3 s 12600 35960 12698 36058 4 gnd
port 3 nsew
rlabel metal3 s 12600 41174 12698 41272 4 gnd
port 3 nsew
rlabel metal3 s 12600 34064 12698 34162 4 gnd
port 3 nsew
rlabel metal3 s 12600 35170 12698 35268 4 gnd
port 3 nsew
rlabel metal3 s 12600 37777 12698 37875 4 gnd
port 3 nsew
rlabel metal3 s 12600 34617 12698 34715 4 gnd
port 3 nsew
rlabel metal3 s 12600 41727 12698 41825 4 gnd
port 3 nsew
rlabel metal3 s 12600 40700 12698 40798 4 gnd
port 3 nsew
rlabel metal3 s 12600 36987 12698 37085 4 gnd
port 3 nsew
rlabel metal3 s 12600 34380 12698 34478 4 gnd
port 3 nsew
rlabel metal3 s 12600 38804 12698 38902 4 gnd
port 3 nsew
rlabel metal3 s 12600 40147 12698 40245 4 gnd
port 3 nsew
rlabel metal3 s 12600 38330 12698 38428 4 gnd
port 3 nsew
rlabel metal3 s 12600 40384 12698 40482 4 gnd
port 3 nsew
rlabel metal3 s 12600 35407 12698 35505 4 gnd
port 3 nsew
rlabel metal3 s 12600 36434 12698 36532 4 gnd
port 3 nsew
rlabel metal3 s 12600 37540 12698 37638 4 gnd
port 3 nsew
rlabel metal3 s 12600 39120 12698 39218 4 gnd
port 3 nsew
rlabel metal3 s 12600 35644 12698 35742 4 gnd
port 3 nsew
rlabel metal3 s 9560 35407 9658 35505 4 gnd
port 3 nsew
rlabel metal3 s 12600 36197 12698 36295 4 gnd
port 3 nsew
rlabel metal3 s 12600 34854 12698 34952 4 gnd
port 3 nsew
rlabel metal3 s 12600 39910 12698 40008 4 gnd
port 3 nsew
rlabel metal3 s 12600 30904 12698 31002 4 gnd
port 3 nsew
rlabel metal3 s 12600 26954 12698 27052 4 gnd
port 3 nsew
rlabel metal3 s 12600 28534 12698 28632 4 gnd
port 3 nsew
rlabel metal3 s 12600 26164 12698 26262 4 gnd
port 3 nsew
rlabel metal3 s 12600 25374 12698 25472 4 gnd
port 3 nsew
rlabel metal3 s 12600 25927 12698 26025 4 gnd
port 3 nsew
rlabel metal3 s 12600 28297 12698 28395 4 gnd
port 3 nsew
rlabel metal3 s 12600 32247 12698 32345 4 gnd
port 3 nsew
rlabel metal3 s 12600 31457 12698 31555 4 gnd
port 3 nsew
rlabel metal3 s 12600 32800 12698 32898 4 gnd
port 3 nsew
rlabel metal3 s 12600 32484 12698 32582 4 gnd
port 3 nsew
rlabel metal3 s 12600 27507 12698 27605 4 gnd
port 3 nsew
rlabel metal3 s 12600 29877 12698 29975 4 gnd
port 3 nsew
rlabel metal3 s 12600 27270 12698 27368 4 gnd
port 3 nsew
rlabel metal3 s 12600 31220 12698 31318 4 gnd
port 3 nsew
rlabel metal3 s 12600 26480 12698 26578 4 gnd
port 3 nsew
rlabel metal3 s 12600 33037 12698 33135 4 gnd
port 3 nsew
rlabel metal3 s 12600 30667 12698 30765 4 gnd
port 3 nsew
rlabel metal3 s 12600 26717 12698 26815 4 gnd
port 3 nsew
rlabel metal3 s 12600 25690 12698 25788 4 gnd
port 3 nsew
rlabel metal3 s 12600 27744 12698 27842 4 gnd
port 3 nsew
rlabel metal3 s 12600 29640 12698 29738 4 gnd
port 3 nsew
rlabel metal3 s 12600 29324 12698 29422 4 gnd
port 3 nsew
rlabel metal3 s 12600 30114 12698 30212 4 gnd
port 3 nsew
rlabel metal3 s 12600 33274 12698 33372 4 gnd
port 3 nsew
rlabel metal3 s 12600 28850 12698 28948 4 gnd
port 3 nsew
rlabel metal3 s 12600 32010 12698 32108 4 gnd
port 3 nsew
rlabel metal3 s 12600 29087 12698 29185 4 gnd
port 3 nsew
rlabel metal3 s 12600 28060 12698 28158 4 gnd
port 3 nsew
rlabel metal3 s 12600 30430 12698 30528 4 gnd
port 3 nsew
rlabel metal3 s 12600 31694 12698 31792 4 gnd
port 3 nsew
rlabel metal3 s 7264 29482 7362 29580 4 gnd
port 3 nsew
rlabel metal3 s 6882 33023 6980 33121 4 vdd
port 2 nsew
rlabel metal3 s 6882 32665 6980 32763 4 vdd
port 2 nsew
rlabel metal3 s 6882 31085 6980 31183 4 vdd
port 2 nsew
rlabel metal3 s 6025 32665 6123 32763 4 gnd
port 3 nsew
rlabel metal3 s 6882 31443 6980 31541 4 vdd
port 2 nsew
rlabel metal3 s 6450 30295 6548 30393 4 vdd
port 2 nsew
rlabel metal3 s 6450 31875 6548 31973 4 vdd
port 2 nsew
rlabel metal3 s 7660 30667 7758 30765 4 vdd
port 2 nsew
rlabel metal3 s 7264 32247 7362 32345 4 gnd
port 3 nsew
rlabel metal3 s 7264 33037 7362 33135 4 gnd
port 3 nsew
rlabel metal3 s 6450 30653 6548 30751 4 vdd
port 2 nsew
rlabel metal3 s 7660 31062 7758 31160 4 vdd
port 2 nsew
rlabel metal3 s 6450 31085 6548 31183 4 vdd
port 2 nsew
rlabel metal3 s 7660 32247 7758 32345 4 vdd
port 2 nsew
rlabel metal3 s 6450 29505 6548 29603 4 vdd
port 2 nsew
rlabel metal3 s 6025 31875 6123 31973 4 gnd
port 3 nsew
rlabel metal3 s 6025 31501 6123 31599 4 gnd
port 3 nsew
rlabel metal3 s 6882 29505 6980 29603 4 vdd
port 2 nsew
rlabel metal3 s 7264 32642 7362 32740 4 gnd
port 3 nsew
rlabel metal3 s 6025 30711 6123 30809 4 gnd
port 3 nsew
rlabel metal3 s 6025 33081 6123 33179 4 gnd
port 3 nsew
rlabel metal3 s 7660 30272 7758 30370 4 vdd
port 2 nsew
rlabel metal3 s 7660 33037 7758 33135 4 vdd
port 2 nsew
rlabel metal3 s 6882 33455 6980 33553 4 vdd
port 2 nsew
rlabel metal3 s 6450 32233 6548 32331 4 vdd
port 2 nsew
rlabel metal3 s 6882 29863 6980 29961 4 vdd
port 2 nsew
rlabel metal3 s 6882 30295 6980 30393 4 vdd
port 2 nsew
rlabel metal3 s 7264 33432 7362 33530 4 gnd
port 3 nsew
rlabel metal3 s 6882 30653 6980 30751 4 vdd
port 2 nsew
rlabel metal3 s 7660 31457 7758 31555 4 vdd
port 2 nsew
rlabel metal3 s 6882 32233 6980 32331 4 vdd
port 2 nsew
rlabel metal3 s 6025 31085 6123 31183 4 gnd
port 3 nsew
rlabel metal3 s 7660 29482 7758 29580 4 vdd
port 2 nsew
rlabel metal3 s 7660 29877 7758 29975 4 vdd
port 2 nsew
rlabel metal3 s 7660 31852 7758 31950 4 vdd
port 2 nsew
rlabel metal3 s 6025 29505 6123 29603 4 gnd
port 3 nsew
rlabel metal3 s 6450 33023 6548 33121 4 vdd
port 2 nsew
rlabel metal3 s 6025 33455 6123 33553 4 gnd
port 3 nsew
rlabel metal3 s 6025 29921 6123 30019 4 gnd
port 3 nsew
rlabel metal3 s 6882 31875 6980 31973 4 vdd
port 2 nsew
rlabel metal3 s 6450 29863 6548 29961 4 vdd
port 2 nsew
rlabel metal3 s 7264 30667 7362 30765 4 gnd
port 3 nsew
rlabel metal3 s 7264 31062 7362 31160 4 gnd
port 3 nsew
rlabel metal3 s 7264 29877 7362 29975 4 gnd
port 3 nsew
rlabel metal3 s 7264 30272 7362 30370 4 gnd
port 3 nsew
rlabel metal3 s 7264 31852 7362 31950 4 gnd
port 3 nsew
rlabel metal3 s 6450 31443 6548 31541 4 vdd
port 2 nsew
rlabel metal3 s 7264 31457 7362 31555 4 gnd
port 3 nsew
rlabel metal3 s 6450 32665 6548 32763 4 vdd
port 2 nsew
rlabel metal3 s 6025 30295 6123 30393 4 gnd
port 3 nsew
rlabel metal3 s 7660 33432 7758 33530 4 vdd
port 2 nsew
rlabel metal3 s 6450 33455 6548 33553 4 vdd
port 2 nsew
rlabel metal3 s 6025 32291 6123 32389 4 gnd
port 3 nsew
rlabel metal3 s 7660 32642 7758 32740 4 vdd
port 2 nsew
rlabel metal3 s 6882 28715 6980 28813 4 vdd
port 2 nsew
rlabel metal3 s 7660 25532 7758 25630 4 vdd
port 2 nsew
rlabel metal3 s 6025 25181 6123 25279 4 gnd
port 3 nsew
rlabel metal3 s 6450 27135 6548 27233 4 vdd
port 2 nsew
rlabel metal3 s 6450 26703 6548 26801 4 vdd
port 2 nsew
rlabel metal3 s 6882 26345 6980 26443 4 vdd
port 2 nsew
rlabel metal3 s 6450 27493 6548 27591 4 vdd
port 2 nsew
rlabel metal3 s 6025 26761 6123 26859 4 gnd
port 3 nsew
rlabel metal3 s 6025 28341 6123 28439 4 gnd
port 3 nsew
rlabel metal3 s 6025 25971 6123 26069 4 gnd
port 3 nsew
rlabel metal3 s 6882 26703 6980 26801 4 vdd
port 2 nsew
rlabel metal3 s 6025 27135 6123 27233 4 gnd
port 3 nsew
rlabel metal3 s 6882 27493 6980 27591 4 vdd
port 2 nsew
rlabel metal3 s 7660 26322 7758 26420 4 vdd
port 2 nsew
rlabel metal3 s 6450 27925 6548 28023 4 vdd
port 2 nsew
rlabel metal3 s 6450 26345 6548 26443 4 vdd
port 2 nsew
rlabel metal3 s 7264 26322 7362 26420 4 gnd
port 3 nsew
rlabel metal3 s 6025 29131 6123 29229 4 gnd
port 3 nsew
rlabel metal3 s 6025 26345 6123 26443 4 gnd
port 3 nsew
rlabel metal3 s 6025 27925 6123 28023 4 gnd
port 3 nsew
rlabel metal3 s 7264 26717 7362 26815 4 gnd
port 3 nsew
rlabel metal3 s 6450 28715 6548 28813 4 vdd
port 2 nsew
rlabel metal3 s 6882 27135 6980 27233 4 vdd
port 2 nsew
rlabel metal3 s 6882 27925 6980 28023 4 vdd
port 2 nsew
rlabel metal3 s 7660 25927 7758 26025 4 vdd
port 2 nsew
rlabel metal3 s 6025 27551 6123 27649 4 gnd
port 3 nsew
rlabel metal3 s 6882 25555 6980 25653 4 vdd
port 2 nsew
rlabel metal3 s 7264 25532 7362 25630 4 gnd
port 3 nsew
rlabel metal3 s 7264 28297 7362 28395 4 gnd
port 3 nsew
rlabel metal3 s 6450 28283 6548 28381 4 vdd
port 2 nsew
rlabel metal3 s 7660 26717 7758 26815 4 vdd
port 2 nsew
rlabel metal3 s 6025 25555 6123 25653 4 gnd
port 3 nsew
rlabel metal3 s 7660 27507 7758 27605 4 vdd
port 2 nsew
rlabel metal3 s 6450 25913 6548 26011 4 vdd
port 2 nsew
rlabel metal3 s 7660 27112 7758 27210 4 vdd
port 2 nsew
rlabel metal3 s 7660 28297 7758 28395 4 vdd
port 2 nsew
rlabel metal3 s 7660 29087 7758 29185 4 vdd
port 2 nsew
rlabel metal3 s 7264 28692 7362 28790 4 gnd
port 3 nsew
rlabel metal3 s 7660 27902 7758 28000 4 vdd
port 2 nsew
rlabel metal3 s 6025 28715 6123 28813 4 gnd
port 3 nsew
rlabel metal3 s 7660 28692 7758 28790 4 vdd
port 2 nsew
rlabel metal3 s 6450 25555 6548 25653 4 vdd
port 2 nsew
rlabel metal3 s 6882 28283 6980 28381 4 vdd
port 2 nsew
rlabel metal3 s 6882 25913 6980 26011 4 vdd
port 2 nsew
rlabel metal3 s 7264 27112 7362 27210 4 gnd
port 3 nsew
rlabel metal3 s 6882 29073 6980 29171 4 vdd
port 2 nsew
rlabel metal3 s 7264 27902 7362 28000 4 gnd
port 3 nsew
rlabel metal3 s 6450 29073 6548 29171 4 vdd
port 2 nsew
rlabel metal3 s 7264 27507 7362 27605 4 gnd
port 3 nsew
rlabel metal3 s 7264 29087 7362 29185 4 gnd
port 3 nsew
rlabel metal3 s 7264 25927 7362 26025 4 gnd
port 3 nsew
rlabel metal3 s 6025 22021 6123 22119 4 gnd
port 3 nsew
rlabel metal3 s 7660 23162 7758 23260 4 vdd
port 2 nsew
rlabel metal3 s 6025 21231 6123 21329 4 gnd
port 3 nsew
rlabel metal3 s 6882 23185 6980 23283 4 vdd
port 2 nsew
rlabel metal3 s 7264 21582 7362 21680 4 gnd
port 3 nsew
rlabel metal3 s 6450 24333 6548 24431 4 vdd
port 2 nsew
rlabel metal3 s 7264 21187 7362 21285 4 gnd
port 3 nsew
rlabel metal3 s 7264 22767 7362 22865 4 gnd
port 3 nsew
rlabel metal3 s 6450 21173 6548 21271 4 vdd
port 2 nsew
rlabel metal3 s 7660 23557 7758 23655 4 vdd
port 2 nsew
rlabel metal3 s 6882 23543 6980 23641 4 vdd
port 2 nsew
rlabel metal3 s 6450 23185 6548 23283 4 vdd
port 2 nsew
rlabel metal3 s 6450 25123 6548 25221 4 vdd
port 2 nsew
rlabel metal3 s 7660 21187 7758 21285 4 vdd
port 2 nsew
rlabel metal3 s 6450 21963 6548 22061 4 vdd
port 2 nsew
rlabel metal3 s 7660 24742 7758 24840 4 vdd
port 2 nsew
rlabel metal3 s 6882 24765 6980 24863 4 vdd
port 2 nsew
rlabel metal3 s 7660 22767 7758 22865 4 vdd
port 2 nsew
rlabel metal3 s 7660 21977 7758 22075 4 vdd
port 2 nsew
rlabel metal3 s 6882 25123 6980 25221 4 vdd
port 2 nsew
rlabel metal3 s 7660 23952 7758 24050 4 vdd
port 2 nsew
rlabel metal3 s 7264 22372 7362 22470 4 gnd
port 3 nsew
rlabel metal3 s 6450 23543 6548 23641 4 vdd
port 2 nsew
rlabel metal3 s 6450 22753 6548 22851 4 vdd
port 2 nsew
rlabel metal3 s 6025 23185 6123 23283 4 gnd
port 3 nsew
rlabel metal3 s 7264 24742 7362 24840 4 gnd
port 3 nsew
rlabel metal3 s 6450 22395 6548 22493 4 vdd
port 2 nsew
rlabel metal3 s 7264 23162 7362 23260 4 gnd
port 3 nsew
rlabel metal3 s 7660 24347 7758 24445 4 vdd
port 2 nsew
rlabel metal3 s 6882 21173 6980 21271 4 vdd
port 2 nsew
rlabel metal3 s 6450 24765 6548 24863 4 vdd
port 2 nsew
rlabel metal3 s 6025 22811 6123 22909 4 gnd
port 3 nsew
rlabel metal3 s 6025 23975 6123 24073 4 gnd
port 3 nsew
rlabel metal3 s 6882 22395 6980 22493 4 vdd
port 2 nsew
rlabel metal3 s 7660 21582 7758 21680 4 vdd
port 2 nsew
rlabel metal3 s 6025 21605 6123 21703 4 gnd
port 3 nsew
rlabel metal3 s 6450 21605 6548 21703 4 vdd
port 2 nsew
rlabel metal3 s 6025 24391 6123 24489 4 gnd
port 3 nsew
rlabel metal3 s 6882 21605 6980 21703 4 vdd
port 2 nsew
rlabel metal3 s 6882 21963 6980 22061 4 vdd
port 2 nsew
rlabel metal3 s 7660 25137 7758 25235 4 vdd
port 2 nsew
rlabel metal3 s 6025 22395 6123 22493 4 gnd
port 3 nsew
rlabel metal3 s 7264 25137 7362 25235 4 gnd
port 3 nsew
rlabel metal3 s 6882 22753 6980 22851 4 vdd
port 2 nsew
rlabel metal3 s 7264 21977 7362 22075 4 gnd
port 3 nsew
rlabel metal3 s 7264 23557 7362 23655 4 gnd
port 3 nsew
rlabel metal3 s 6882 23975 6980 24073 4 vdd
port 2 nsew
rlabel metal3 s 7264 23952 7362 24050 4 gnd
port 3 nsew
rlabel metal3 s 7264 24347 7362 24445 4 gnd
port 3 nsew
rlabel metal3 s 6025 24765 6123 24863 4 gnd
port 3 nsew
rlabel metal3 s 6450 23975 6548 24073 4 vdd
port 2 nsew
rlabel metal3 s 7660 22372 7758 22470 4 vdd
port 2 nsew
rlabel metal3 s 6882 24333 6980 24431 4 vdd
port 2 nsew
rlabel metal3 s 6025 23601 6123 23699 4 gnd
port 3 nsew
rlabel metal3 s 2611 16865 2709 16963 4 gnd
port 3 nsew
rlabel metal3 s 4246 17632 4344 17730 4 vdd
port 2 nsew
rlabel metal3 s 3468 16865 3566 16963 4 vdd
port 2 nsew
rlabel metal3 s 3850 16842 3948 16940 4 gnd
port 3 nsew
rlabel metal3 s 3036 16865 3134 16963 4 vdd
port 2 nsew
rlabel metal3 s 2611 17655 2709 17753 4 gnd
port 3 nsew
rlabel metal3 s 3468 17655 3566 17753 4 vdd
port 2 nsew
rlabel metal3 s 4246 16842 4344 16940 4 vdd
port 2 nsew
rlabel metal3 s 3850 17632 3948 17730 4 gnd
port 3 nsew
rlabel metal3 s 3036 17655 3134 17753 4 vdd
port 2 nsew
rlabel metal3 s 6450 16865 6548 16963 4 vdd
port 2 nsew
rlabel metal3 s 7660 19607 7758 19705 4 vdd
port 2 nsew
rlabel metal3 s 6450 17223 6548 17321 4 vdd
port 2 nsew
rlabel metal3 s 6882 18803 6980 18901 4 vdd
port 2 nsew
rlabel metal3 s 6025 18445 6123 18543 4 gnd
port 3 nsew
rlabel metal3 s 6882 20025 6980 20123 4 vdd
port 2 nsew
rlabel metal3 s 6450 18013 6548 18111 4 vdd
port 2 nsew
rlabel metal3 s 6882 20383 6980 20481 4 vdd
port 2 nsew
rlabel metal3 s 6450 18445 6548 18543 4 vdd
port 2 nsew
rlabel metal3 s 7264 16842 7362 16940 4 gnd
port 3 nsew
rlabel metal3 s 7264 18422 7362 18520 4 gnd
port 3 nsew
rlabel metal3 s 6450 20383 6548 20481 4 vdd
port 2 nsew
rlabel metal3 s 7264 20397 7362 20495 4 gnd
port 3 nsew
rlabel metal3 s 7660 19212 7758 19310 4 vdd
port 2 nsew
rlabel metal3 s 7660 20002 7758 20100 4 vdd
port 2 nsew
rlabel metal3 s 6025 19651 6123 19749 4 gnd
port 3 nsew
rlabel metal3 s 7660 17237 7758 17335 4 vdd
port 2 nsew
rlabel metal3 s 6882 19235 6980 19333 4 vdd
port 2 nsew
rlabel metal3 s 6450 18803 6548 18901 4 vdd
port 2 nsew
rlabel metal3 s 7660 17632 7758 17730 4 vdd
port 2 nsew
rlabel metal3 s 6882 17655 6980 17753 4 vdd
port 2 nsew
rlabel metal3 s 6450 19235 6548 19333 4 vdd
port 2 nsew
rlabel metal3 s 6882 20815 6980 20913 4 vdd
port 2 nsew
rlabel metal3 s 7660 18817 7758 18915 4 vdd
port 2 nsew
rlabel metal3 s 6025 16865 6123 16963 4 gnd
port 3 nsew
rlabel metal3 s 6025 20025 6123 20123 4 gnd
port 3 nsew
rlabel metal3 s 6882 17223 6980 17321 4 vdd
port 2 nsew
rlabel metal3 s 6450 20025 6548 20123 4 vdd
port 2 nsew
rlabel metal3 s 7264 19212 7362 19310 4 gnd
port 3 nsew
rlabel metal3 s 7660 18422 7758 18520 4 vdd
port 2 nsew
rlabel metal3 s 6450 19593 6548 19691 4 vdd
port 2 nsew
rlabel metal3 s 6025 17655 6123 17753 4 gnd
port 3 nsew
rlabel metal3 s 6025 18071 6123 18169 4 gnd
port 3 nsew
rlabel metal3 s 6882 18013 6980 18111 4 vdd
port 2 nsew
rlabel metal3 s 6882 18445 6980 18543 4 vdd
port 2 nsew
rlabel metal3 s 7660 16842 7758 16940 4 vdd
port 2 nsew
rlabel metal3 s 6450 20815 6548 20913 4 vdd
port 2 nsew
rlabel metal3 s 6025 17281 6123 17379 4 gnd
port 3 nsew
rlabel metal3 s 6025 20441 6123 20539 4 gnd
port 3 nsew
rlabel metal3 s 7264 18027 7362 18125 4 gnd
port 3 nsew
rlabel metal3 s 7660 20397 7758 20495 4 vdd
port 2 nsew
rlabel metal3 s 7660 18027 7758 18125 4 vdd
port 2 nsew
rlabel metal3 s 6025 20815 6123 20913 4 gnd
port 3 nsew
rlabel metal3 s 6882 19593 6980 19691 4 vdd
port 2 nsew
rlabel metal3 s 6882 16865 6980 16963 4 vdd
port 2 nsew
rlabel metal3 s 7264 19607 7362 19705 4 gnd
port 3 nsew
rlabel metal3 s 7264 17632 7362 17730 4 gnd
port 3 nsew
rlabel metal3 s 7264 20792 7362 20890 4 gnd
port 3 nsew
rlabel metal3 s 7660 20792 7758 20890 4 vdd
port 2 nsew
rlabel metal3 s 6025 18861 6123 18959 4 gnd
port 3 nsew
rlabel metal3 s 6025 19235 6123 19333 4 gnd
port 3 nsew
rlabel metal3 s 7264 20002 7362 20100 4 gnd
port 3 nsew
rlabel metal3 s 7264 18817 7362 18915 4 gnd
port 3 nsew
rlabel metal3 s 7264 17237 7362 17335 4 gnd
port 3 nsew
rlabel metal3 s 6450 17655 6548 17753 4 vdd
port 2 nsew
rlabel metal3 s 12600 20397 12698 20495 4 gnd
port 3 nsew
rlabel metal3 s 12600 22767 12698 22865 4 gnd
port 3 nsew
rlabel metal3 s 12600 17237 12698 17335 4 gnd
port 3 nsew
rlabel metal3 s 12600 18264 12698 18362 4 gnd
port 3 nsew
rlabel metal3 s 12600 20950 12698 21048 4 gnd
port 3 nsew
rlabel metal3 s 12600 22530 12698 22628 4 gnd
port 3 nsew
rlabel metal3 s 12600 24900 12698 24998 4 gnd
port 3 nsew
rlabel metal3 s 12600 24347 12698 24445 4 gnd
port 3 nsew
rlabel metal3 s 12600 21740 12698 21838 4 gnd
port 3 nsew
rlabel metal3 s 12600 17790 12698 17888 4 gnd
port 3 nsew
rlabel metal3 s 12600 21424 12698 21522 4 gnd
port 3 nsew
rlabel metal3 s 12600 24584 12698 24682 4 gnd
port 3 nsew
rlabel metal3 s 12600 24110 12698 24208 4 gnd
port 3 nsew
rlabel metal3 s 12600 18580 12698 18678 4 gnd
port 3 nsew
rlabel metal3 s 12600 21187 12698 21285 4 gnd
port 3 nsew
rlabel metal3 s 12600 20160 12698 20258 4 gnd
port 3 nsew
rlabel metal3 s 12600 19844 12698 19942 4 gnd
port 3 nsew
rlabel metal3 s 12600 23794 12698 23892 4 gnd
port 3 nsew
rlabel metal3 s 12600 23004 12698 23102 4 gnd
port 3 nsew
rlabel metal3 s 12600 19054 12698 19152 4 gnd
port 3 nsew
rlabel metal3 s 12600 18817 12698 18915 4 gnd
port 3 nsew
rlabel metal3 s 12600 21977 12698 22075 4 gnd
port 3 nsew
rlabel metal3 s 12600 19607 12698 19705 4 gnd
port 3 nsew
rlabel metal3 s 12600 20634 12698 20732 4 gnd
port 3 nsew
rlabel metal3 s 12600 25137 12698 25235 4 gnd
port 3 nsew
rlabel metal3 s 12600 17474 12698 17572 4 gnd
port 3 nsew
rlabel metal3 s 12600 18027 12698 18125 4 gnd
port 3 nsew
rlabel metal3 s 12600 19370 12698 19468 4 gnd
port 3 nsew
rlabel metal3 s 12600 22214 12698 22312 4 gnd
port 3 nsew
rlabel metal3 s 12600 23320 12698 23418 4 gnd
port 3 nsew
rlabel metal3 s 12600 23557 12698 23655 4 gnd
port 3 nsew
rlabel metal3 s 12600 17000 12698 17098 4 gnd
port 3 nsew
rlabel metal3 s 15168 9566 15266 9664 4 vdd
port 2 nsew
rlabel metal3 s 15911 8975 16009 9073 4 vdd
port 2 nsew
rlabel metal3 s 15792 9566 15890 9664 4 vdd
port 2 nsew
rlabel metal3 s 14663 8975 14761 9073 4 vdd
port 2 nsew
rlabel metal3 s 12600 13524 12698 13622 4 gnd
port 3 nsew
rlabel metal3 s 17040 9566 17138 9664 4 vdd
port 2 nsew
rlabel metal3 s 12600 15104 12698 15202 4 gnd
port 3 nsew
rlabel metal3 s 12600 15894 12698 15992 4 gnd
port 3 nsew
rlabel metal3 s 12600 14867 12698 14965 4 gnd
port 3 nsew
rlabel metal3 s 12600 16210 12698 16308 4 gnd
port 3 nsew
rlabel metal3 s 12600 12260 12698 12358 4 gnd
port 3 nsew
rlabel metal3 s 12234 10000 12332 10098 4 gnd
port 3 nsew
rlabel metal3 s 13801 8975 13899 9073 4 vdd
port 2 nsew
rlabel metal3 s 17159 8975 17257 9073 4 vdd
port 2 nsew
rlabel metal3 s 12600 16447 12698 16545 4 gnd
port 3 nsew
rlabel metal3 s 12600 15657 12698 15755 4 gnd
port 3 nsew
rlabel metal3 s 11208 9930 11306 10028 4 vdd
port 2 nsew
rlabel metal3 s 14544 9566 14642 9664 4 vdd
port 2 nsew
rlabel metal3 s 13415 8975 13513 9073 4 vdd
port 2 nsew
rlabel metal3 s 16416 9566 16514 9664 4 vdd
port 2 nsew
rlabel metal3 s 13920 9566 14018 9664 4 vdd
port 2 nsew
rlabel metal3 s 12600 10917 12698 11015 4 gnd
port 3 nsew
rlabel metal3 s 12600 15420 12698 15518 4 gnd
port 3 nsew
rlabel metal3 s 16297 8975 16395 9073 4 vdd
port 2 nsew
rlabel metal3 s 12600 11470 12698 11568 4 gnd
port 3 nsew
rlabel metal3 s 12600 11154 12698 11252 4 gnd
port 3 nsew
rlabel metal3 s 12600 12734 12698 12832 4 gnd
port 3 nsew
rlabel metal3 s 12600 14314 12698 14412 4 gnd
port 3 nsew
rlabel metal3 s 12600 12497 12698 12595 4 gnd
port 3 nsew
rlabel metal3 s 12600 10127 12698 10225 4 gnd
port 3 nsew
rlabel metal3 s 12600 13050 12698 13148 4 gnd
port 3 nsew
rlabel metal3 s 12600 13287 12698 13385 4 gnd
port 3 nsew
rlabel metal3 s 12600 16684 12698 16782 4 gnd
port 3 nsew
rlabel metal3 s 13296 9566 13394 9664 4 vdd
port 2 nsew
rlabel metal3 s 12600 13840 12698 13938 4 gnd
port 3 nsew
rlabel metal3 s 12600 10364 12698 10462 4 gnd
port 3 nsew
rlabel metal3 s 15049 8975 15147 9073 4 vdd
port 2 nsew
rlabel metal3 s 12600 11944 12698 12042 4 gnd
port 3 nsew
rlabel metal3 s 12600 14630 12698 14728 4 gnd
port 3 nsew
rlabel metal3 s 12600 14077 12698 14175 4 gnd
port 3 nsew
rlabel metal3 s 12600 11707 12698 11805 4 gnd
port 3 nsew
rlabel metal3 s 12600 10680 12698 10778 4 gnd
port 3 nsew
rlabel metal3 s 7264 14472 7362 14570 4 gnd
port 3 nsew
rlabel metal3 s 7264 13287 7362 13385 4 gnd
port 3 nsew
rlabel metal3 s 6025 12915 6123 13013 4 gnd
port 3 nsew
rlabel metal3 s 6025 16491 6123 16589 4 gnd
port 3 nsew
rlabel metal3 s 6450 13273 6548 13371 4 vdd
port 2 nsew
rlabel metal3 s 6450 16075 6548 16173 4 vdd
port 2 nsew
rlabel metal3 s 6882 13273 6980 13371 4 vdd
port 2 nsew
rlabel metal3 s 7264 15657 7362 15755 4 gnd
port 3 nsew
rlabel metal3 s 6882 14495 6980 14593 4 vdd
port 2 nsew
rlabel metal3 s 6025 13331 6123 13429 4 gnd
port 3 nsew
rlabel metal3 s 6025 16075 6123 16173 4 gnd
port 3 nsew
rlabel metal3 s 6882 15643 6980 15741 4 vdd
port 2 nsew
rlabel metal3 s 6882 16433 6980 16531 4 vdd
port 2 nsew
rlabel metal3 s 7660 13682 7758 13780 4 vdd
port 2 nsew
rlabel metal3 s 6025 15701 6123 15799 4 gnd
port 3 nsew
rlabel metal3 s 7660 14077 7758 14175 4 vdd
port 2 nsew
rlabel metal3 s 6025 14121 6123 14219 4 gnd
port 3 nsew
rlabel metal3 s 6450 15285 6548 15383 4 vdd
port 2 nsew
rlabel metal3 s 6882 13705 6980 13803 4 vdd
port 2 nsew
rlabel metal3 s 6025 14911 6123 15009 4 gnd
port 3 nsew
rlabel metal3 s 7660 14867 7758 14965 4 vdd
port 2 nsew
rlabel metal3 s 6882 16075 6980 16173 4 vdd
port 2 nsew
rlabel metal3 s 7660 15657 7758 15755 4 vdd
port 2 nsew
rlabel metal3 s 6882 14063 6980 14161 4 vdd
port 2 nsew
rlabel metal3 s 7660 16447 7758 16545 4 vdd
port 2 nsew
rlabel metal3 s 6882 14853 6980 14951 4 vdd
port 2 nsew
rlabel metal3 s 6025 13705 6123 13803 4 gnd
port 3 nsew
rlabel metal3 s 7264 14077 7362 14175 4 gnd
port 3 nsew
rlabel metal3 s 6882 12915 6980 13013 4 vdd
port 2 nsew
rlabel metal3 s 6882 15285 6980 15383 4 vdd
port 2 nsew
rlabel metal3 s 7264 16052 7362 16150 4 gnd
port 3 nsew
rlabel metal3 s 6450 14495 6548 14593 4 vdd
port 2 nsew
rlabel metal3 s 7660 13287 7758 13385 4 vdd
port 2 nsew
rlabel metal3 s 6450 12915 6548 13013 4 vdd
port 2 nsew
rlabel metal3 s 6450 13705 6548 13803 4 vdd
port 2 nsew
rlabel metal3 s 6025 14495 6123 14593 4 gnd
port 3 nsew
rlabel metal3 s 7264 15262 7362 15360 4 gnd
port 3 nsew
rlabel metal3 s 6025 15285 6123 15383 4 gnd
port 3 nsew
rlabel metal3 s 6450 14063 6548 14161 4 vdd
port 2 nsew
rlabel metal3 s 6450 15643 6548 15741 4 vdd
port 2 nsew
rlabel metal3 s 6450 14853 6548 14951 4 vdd
port 2 nsew
rlabel metal3 s 7264 14867 7362 14965 4 gnd
port 3 nsew
rlabel metal3 s 7660 16052 7758 16150 4 vdd
port 2 nsew
rlabel metal3 s 7660 12892 7758 12990 4 vdd
port 2 nsew
rlabel metal3 s 7660 14472 7758 14570 4 vdd
port 2 nsew
rlabel metal3 s 6450 16433 6548 16531 4 vdd
port 2 nsew
rlabel metal3 s 7264 12892 7362 12990 4 gnd
port 3 nsew
rlabel metal3 s 7264 16447 7362 16545 4 gnd
port 3 nsew
rlabel metal3 s 7660 15262 7758 15360 4 vdd
port 2 nsew
rlabel metal3 s 7264 13682 7362 13780 4 gnd
port 3 nsew
rlabel metal3 s 1752 12892 1850 12990 4 gnd
port 3 nsew
rlabel metal3 s 2148 12892 2246 12990 4 vdd
port 2 nsew
rlabel metal3 s 2611 16075 2709 16173 4 gnd
port 3 nsew
rlabel metal3 s 3468 16075 3566 16173 4 vdd
port 2 nsew
rlabel metal3 s 3046 12899 3144 12997 4 gnd
port 3 nsew
rlabel metal3 s 3850 13682 3948 13780 4 gnd
port 3 nsew
rlabel metal3 s 3046 13689 3144 13787 4 gnd
port 3 nsew
rlabel metal3 s 4246 13682 4344 13780 4 vdd
port 2 nsew
rlabel metal3 s 4246 15262 4344 15360 4 vdd
port 2 nsew
rlabel metal3 s 3468 15285 3566 15383 4 vdd
port 2 nsew
rlabel metal3 s 3850 12892 3948 12990 4 gnd
port 3 nsew
rlabel metal3 s 3471 12899 3569 12997 4 vdd
port 2 nsew
rlabel metal3 s 3471 13689 3569 13787 4 vdd
port 2 nsew
rlabel metal3 s 4246 16052 4344 16150 4 vdd
port 2 nsew
rlabel metal3 s 4246 12892 4344 12990 4 vdd
port 2 nsew
rlabel metal3 s 1156 15262 1254 15360 4 gnd
port 3 nsew
rlabel metal3 s 2611 15285 2709 15383 4 gnd
port 3 nsew
rlabel metal3 s 3850 15262 3948 15360 4 gnd
port 3 nsew
rlabel metal3 s 1552 15262 1650 15360 4 vdd
port 2 nsew
rlabel metal3 s 3036 15285 3134 15383 4 vdd
port 2 nsew
rlabel metal3 s 3850 16052 3948 16150 4 gnd
port 3 nsew
rlabel metal3 s 3036 16075 3134 16173 4 vdd
port 2 nsew
rlabel metal3 s 3850 11312 3948 11410 4 gnd
port 3 nsew
rlabel metal3 s 3046 11319 3144 11417 4 gnd
port 3 nsew
rlabel metal3 s 3046 10529 3144 10627 4 gnd
port 3 nsew
rlabel metal3 s 2148 10522 2246 10620 4 vdd
port 2 nsew
rlabel metal3 s 1752 10522 1850 10620 4 gnd
port 3 nsew
rlabel metal3 s 4246 10522 4344 10620 4 vdd
port 2 nsew
rlabel metal3 s 3471 11319 3569 11417 4 vdd
port 2 nsew
rlabel metal3 s 4246 11312 4344 11410 4 vdd
port 2 nsew
rlabel metal3 s 3471 10529 3569 10627 4 vdd
port 2 nsew
rlabel metal3 s 3850 10522 3948 10620 4 gnd
port 3 nsew
rlabel metal3 s 6025 12125 6123 12223 4 gnd
port 3 nsew
rlabel metal3 s 6025 12541 6123 12639 4 gnd
port 3 nsew
rlabel metal3 s 6450 10903 6548 11001 4 vdd
port 2 nsew
rlabel metal3 s 6882 10903 6980 11001 4 vdd
port 2 nsew
rlabel metal3 s 7660 11312 7758 11410 4 vdd
port 2 nsew
rlabel metal3 s 6882 10545 6980 10643 4 vdd
port 2 nsew
rlabel metal3 s 7264 12497 7362 12595 4 gnd
port 3 nsew
rlabel metal3 s 7264 12102 7362 12200 4 gnd
port 3 nsew
rlabel metal3 s 6025 11335 6123 11433 4 gnd
port 3 nsew
rlabel metal3 s 6450 12125 6548 12223 4 vdd
port 2 nsew
rlabel metal3 s 7660 12497 7758 12595 4 vdd
port 2 nsew
rlabel metal3 s 6450 11335 6548 11433 4 vdd
port 2 nsew
rlabel metal3 s 6882 12125 6980 12223 4 vdd
port 2 nsew
rlabel metal3 s 6025 11751 6123 11849 4 gnd
port 3 nsew
rlabel metal3 s 6450 11693 6548 11791 4 vdd
port 2 nsew
rlabel metal3 s 7264 11312 7362 11410 4 gnd
port 3 nsew
rlabel metal3 s 7264 11707 7362 11805 4 gnd
port 3 nsew
rlabel metal3 s 6025 10961 6123 11059 4 gnd
port 3 nsew
rlabel metal3 s 7660 10522 7758 10620 4 vdd
port 2 nsew
rlabel metal3 s 6450 10545 6548 10643 4 vdd
port 2 nsew
rlabel metal3 s 7685 9936 7783 10034 4 vdd
port 2 nsew
rlabel metal3 s 6450 12483 6548 12581 4 vdd
port 2 nsew
rlabel metal3 s 7264 10917 7362 11015 4 gnd
port 3 nsew
rlabel metal3 s 7264 10522 7362 10620 4 gnd
port 3 nsew
rlabel metal3 s 8517 9942 8615 10040 4 vdd
port 2 nsew
rlabel metal3 s 6882 12483 6980 12581 4 vdd
port 2 nsew
rlabel metal3 s 6882 11693 6980 11791 4 vdd
port 2 nsew
rlabel metal3 s 7660 11707 7758 11805 4 vdd
port 2 nsew
rlabel metal3 s 6025 10545 6123 10643 4 gnd
port 3 nsew
rlabel metal3 s 7660 10917 7758 11015 4 vdd
port 2 nsew
rlabel metal3 s 7660 12102 7758 12200 4 vdd
port 2 nsew
rlabel metal3 s 6882 11335 6980 11433 4 vdd
port 2 nsew
rlabel metal3 s 6708 4758 6806 4856 4 gnd
port 3 nsew
rlabel metal3 s 0 8226 13577 8286 4 rbl_bl_0_0
port 4 nsew
rlabel metal3 s 6708 6172 6806 6270 4 vdd
port 2 nsew
rlabel metal3 s 6708 7586 6806 7684 4 gnd
port 3 nsew
rlabel metal3 s 16366 1979 16464 2077 4 gnd
port 3 nsew
rlabel metal3 s 12234 1120 12332 1218 4 vdd
port 2 nsew
rlabel metal3 s 13977 4903 14075 5001 4 vdd
port 2 nsew
rlabel metal3 s 13989 3743 14087 3841 4 gnd
port 3 nsew
rlabel metal3 s 13884 1563 13982 1661 4 vdd
port 2 nsew
rlabel metal3 s 16485 3743 16583 3841 4 gnd
port 3 nsew
rlabel metal3 s 13864 2513 13962 2611 4 vdd
port 2 nsew
rlabel metal3 s 14059 5677 14157 5775 4 gnd
port 3 nsew
rlabel metal3 s 15237 3743 15335 3841 4 gnd
port 3 nsew
rlabel metal3 s 15225 4903 15323 5001 4 vdd
port 2 nsew
rlabel metal3 s 16371 2950 16469 3048 4 gnd
port 3 nsew
rlabel metal3 s 14232 7426 14330 7524 4 gnd
port 3 nsew
rlabel metal3 s 12234 0 12332 98 4 gnd
port 3 nsew
rlabel metal3 s 16380 1563 16478 1661 4 vdd
port 2 nsew
rlabel metal3 s 16485 4065 16583 4163 4 vdd
port 2 nsew
rlabel metal3 s 16473 4903 16571 5001 4 vdd
port 2 nsew
rlabel metal3 s 13989 4065 14087 4163 4 vdd
port 2 nsew
rlabel metal3 s 13875 2950 13973 3048 4 gnd
port 3 nsew
rlabel metal3 s 15118 1979 15216 2077 4 gnd
port 3 nsew
rlabel metal3 s 15480 7426 15578 7524 4 gnd
port 3 nsew
rlabel metal3 s 16481 2181 16579 2279 4 gnd
port 3 nsew
rlabel metal3 s 15307 5677 15405 5775 4 gnd
port 3 nsew
rlabel metal3 s 13870 1979 13968 2077 4 gnd
port 3 nsew
rlabel metal3 s 16360 2513 16458 2611 4 vdd
port 2 nsew
rlabel metal3 s 13985 2181 14083 2279 4 gnd
port 3 nsew
rlabel metal3 s 16555 5677 16653 5775 4 gnd
port 3 nsew
rlabel metal3 s 15233 2181 15331 2279 4 gnd
port 3 nsew
rlabel metal3 s 15132 1563 15230 1661 4 vdd
port 2 nsew
rlabel metal3 s 15237 4065 15335 4163 4 vdd
port 2 nsew
rlabel metal3 s 15123 2950 15221 3048 4 gnd
port 3 nsew
rlabel metal3 s 16728 7426 16826 7524 4 gnd
port 3 nsew
rlabel metal3 s 15112 2513 15210 2611 4 vdd
port 2 nsew
rlabel metal3 s 25895 8975 25993 9073 4 vdd
port 2 nsew
rlabel metal3 s 27648 9566 27746 9664 4 vdd
port 2 nsew
rlabel metal3 s 31273 8975 31371 9073 4 vdd
port 2 nsew
rlabel metal3 s 29520 9566 29618 9664 4 vdd
port 2 nsew
rlabel metal3 s 27024 9566 27122 9664 4 vdd
port 2 nsew
rlabel metal3 s 32135 8975 32233 9073 4 vdd
port 2 nsew
rlabel metal3 s 33383 8975 33481 9073 4 vdd
port 2 nsew
rlabel metal3 s 28896 9566 28994 9664 4 vdd
port 2 nsew
rlabel metal3 s 26400 9566 26498 9664 4 vdd
port 2 nsew
rlabel metal3 s 28391 8975 28489 9073 4 vdd
port 2 nsew
rlabel metal3 s 30144 9566 30242 9664 4 vdd
port 2 nsew
rlabel metal3 s 26281 8975 26379 9073 4 vdd
port 2 nsew
rlabel metal3 s 32521 8975 32619 9073 4 vdd
port 2 nsew
rlabel metal3 s 27143 8975 27241 9073 4 vdd
port 2 nsew
rlabel metal3 s 33264 9566 33362 9664 4 vdd
port 2 nsew
rlabel metal3 s 30887 8975 30985 9073 4 vdd
port 2 nsew
rlabel metal3 s 31392 9566 31490 9664 4 vdd
port 2 nsew
rlabel metal3 s 32016 9566 32114 9664 4 vdd
port 2 nsew
rlabel metal3 s 28777 8975 28875 9073 4 vdd
port 2 nsew
rlabel metal3 s 28272 9566 28370 9664 4 vdd
port 2 nsew
rlabel metal3 s 32640 9566 32738 9664 4 vdd
port 2 nsew
rlabel metal3 s 30025 8975 30123 9073 4 vdd
port 2 nsew
rlabel metal3 s 27529 8975 27627 9073 4 vdd
port 2 nsew
rlabel metal3 s 29639 8975 29737 9073 4 vdd
port 2 nsew
rlabel metal3 s 30768 9566 30866 9664 4 vdd
port 2 nsew
rlabel metal3 s 25776 9566 25874 9664 4 vdd
port 2 nsew
rlabel metal3 s 20041 8975 20139 9073 4 vdd
port 2 nsew
rlabel metal3 s 23904 9566 24002 9664 4 vdd
port 2 nsew
rlabel metal3 s 17545 8975 17643 9073 4 vdd
port 2 nsew
rlabel metal3 s 25152 9566 25250 9664 4 vdd
port 2 nsew
rlabel metal3 s 20160 9566 20258 9664 4 vdd
port 2 nsew
rlabel metal3 s 18407 8975 18505 9073 4 vdd
port 2 nsew
rlabel metal3 s 22151 8975 22249 9073 4 vdd
port 2 nsew
rlabel metal3 s 21289 8975 21387 9073 4 vdd
port 2 nsew
rlabel metal3 s 22656 9566 22754 9664 4 vdd
port 2 nsew
rlabel metal3 s 23399 8975 23497 9073 4 vdd
port 2 nsew
rlabel metal3 s 24528 9566 24626 9664 4 vdd
port 2 nsew
rlabel metal3 s 19536 9566 19634 9664 4 vdd
port 2 nsew
rlabel metal3 s 25033 8975 25131 9073 4 vdd
port 2 nsew
rlabel metal3 s 22537 8975 22635 9073 4 vdd
port 2 nsew
rlabel metal3 s 20903 8975 21001 9073 4 vdd
port 2 nsew
rlabel metal3 s 18793 8975 18891 9073 4 vdd
port 2 nsew
rlabel metal3 s 22032 9566 22130 9664 4 vdd
port 2 nsew
rlabel metal3 s 20784 9566 20882 9664 4 vdd
port 2 nsew
rlabel metal3 s 24647 8975 24745 9073 4 vdd
port 2 nsew
rlabel metal3 s 17664 9566 17762 9664 4 vdd
port 2 nsew
rlabel metal3 s 21408 9566 21506 9664 4 vdd
port 2 nsew
rlabel metal3 s 23280 9566 23378 9664 4 vdd
port 2 nsew
rlabel metal3 s 23785 8975 23883 9073 4 vdd
port 2 nsew
rlabel metal3 s 19655 8975 19753 9073 4 vdd
port 2 nsew
rlabel metal3 s 18912 9566 19010 9664 4 vdd
port 2 nsew
rlabel metal3 s 18288 9566 18386 9664 4 vdd
port 2 nsew
rlabel metal3 s 18981 4065 19079 4163 4 vdd
port 2 nsew
rlabel metal3 s 17628 1563 17726 1661 4 vdd
port 2 nsew
rlabel metal3 s 22611 2950 22709 3048 4 gnd
port 3 nsew
rlabel metal3 s 23973 4065 24071 4163 4 vdd
port 2 nsew
rlabel metal3 s 17803 5677 17901 5775 4 gnd
port 3 nsew
rlabel metal3 s 25221 4065 25319 4163 4 vdd
port 2 nsew
rlabel metal3 s 25096 2513 25194 2611 4 vdd
port 2 nsew
rlabel metal3 s 23854 1979 23952 2077 4 gnd
port 3 nsew
rlabel metal3 s 19224 7426 19322 7524 4 gnd
port 3 nsew
rlabel metal3 s 20299 5677 20397 5775 4 gnd
port 3 nsew
rlabel metal3 s 20115 2950 20213 3048 4 gnd
port 3 nsew
rlabel metal3 s 25217 2181 25315 2279 4 gnd
port 3 nsew
rlabel metal3 s 20229 3743 20327 3841 4 gnd
port 3 nsew
rlabel metal3 s 18969 4903 19067 5001 4 vdd
port 2 nsew
rlabel metal3 s 23969 2181 24067 2279 4 gnd
port 3 nsew
rlabel metal3 s 17608 2513 17706 2611 4 vdd
port 2 nsew
rlabel metal3 s 17733 3743 17831 3841 4 gnd
port 3 nsew
rlabel metal3 s 25107 2950 25205 3048 4 gnd
port 3 nsew
rlabel metal3 s 18876 1563 18974 1661 4 vdd
port 2 nsew
rlabel metal3 s 21477 3743 21575 3841 4 gnd
port 3 nsew
rlabel metal3 s 21465 4903 21563 5001 4 vdd
port 2 nsew
rlabel metal3 s 25291 5677 25389 5775 4 gnd
port 3 nsew
rlabel metal3 s 20217 4903 20315 5001 4 vdd
port 2 nsew
rlabel metal3 s 25209 4903 25307 5001 4 vdd
port 2 nsew
rlabel metal3 s 20225 2181 20323 2279 4 gnd
port 3 nsew
rlabel metal3 s 24216 7426 24314 7524 4 gnd
port 3 nsew
rlabel metal3 s 21372 1563 21470 1661 4 vdd
port 2 nsew
rlabel metal3 s 18977 2181 19075 2279 4 gnd
port 3 nsew
rlabel metal3 s 25102 1979 25200 2077 4 gnd
port 3 nsew
rlabel metal3 s 20472 7426 20570 7524 4 gnd
port 3 nsew
rlabel metal3 s 22713 4903 22811 5001 4 vdd
port 2 nsew
rlabel metal3 s 20110 1979 20208 2077 4 gnd
port 3 nsew
rlabel metal3 s 18862 1979 18960 2077 4 gnd
port 3 nsew
rlabel metal3 s 21358 1979 21456 2077 4 gnd
port 3 nsew
rlabel metal3 s 18856 2513 18954 2611 4 vdd
port 2 nsew
rlabel metal3 s 25116 1563 25214 1661 4 vdd
port 2 nsew
rlabel metal3 s 18981 3743 19079 3841 4 gnd
port 3 nsew
rlabel metal3 s 22725 4065 22823 4163 4 vdd
port 2 nsew
rlabel metal3 s 25221 3743 25319 3841 4 gnd
port 3 nsew
rlabel metal3 s 24043 5677 24141 5775 4 gnd
port 3 nsew
rlabel metal3 s 21473 2181 21571 2279 4 gnd
port 3 nsew
rlabel metal3 s 23973 3743 24071 3841 4 gnd
port 3 nsew
rlabel metal3 s 17619 2950 17717 3048 4 gnd
port 3 nsew
rlabel metal3 s 22606 1979 22704 2077 4 gnd
port 3 nsew
rlabel metal3 s 25464 7426 25562 7524 4 gnd
port 3 nsew
rlabel metal3 s 17733 4065 17831 4163 4 vdd
port 2 nsew
rlabel metal3 s 20124 1563 20222 1661 4 vdd
port 2 nsew
rlabel metal3 s 21720 7426 21818 7524 4 gnd
port 3 nsew
rlabel metal3 s 22600 2513 22698 2611 4 vdd
port 2 nsew
rlabel metal3 s 22968 7426 23066 7524 4 gnd
port 3 nsew
rlabel metal3 s 17614 1979 17712 2077 4 gnd
port 3 nsew
rlabel metal3 s 17976 7426 18074 7524 4 gnd
port 3 nsew
rlabel metal3 s 22721 2181 22819 2279 4 gnd
port 3 nsew
rlabel metal3 s 17729 2181 17827 2279 4 gnd
port 3 nsew
rlabel metal3 s 22725 3743 22823 3841 4 gnd
port 3 nsew
rlabel metal3 s 23848 2513 23946 2611 4 vdd
port 2 nsew
rlabel metal3 s 23961 4903 24059 5001 4 vdd
port 2 nsew
rlabel metal3 s 21477 4065 21575 4163 4 vdd
port 2 nsew
rlabel metal3 s 20229 4065 20327 4163 4 vdd
port 2 nsew
rlabel metal3 s 22620 1563 22718 1661 4 vdd
port 2 nsew
rlabel metal3 s 23868 1563 23966 1661 4 vdd
port 2 nsew
rlabel metal3 s 22795 5677 22893 5775 4 gnd
port 3 nsew
rlabel metal3 s 18867 2950 18965 3048 4 gnd
port 3 nsew
rlabel metal3 s 21352 2513 21450 2611 4 vdd
port 2 nsew
rlabel metal3 s 20104 2513 20202 2611 4 vdd
port 2 nsew
rlabel metal3 s 19051 5677 19149 5775 4 gnd
port 3 nsew
rlabel metal3 s 23859 2950 23957 3048 4 gnd
port 3 nsew
rlabel metal3 s 21547 5677 21645 5775 4 gnd
port 3 nsew
rlabel metal3 s 21363 2950 21461 3048 4 gnd
port 3 nsew
rlabel metal3 s 17721 4903 17819 5001 4 vdd
port 2 nsew
rlabel metal3 s 26469 3743 26567 3841 4 gnd
port 3 nsew
rlabel metal3 s 27612 1563 27710 1661 4 vdd
port 2 nsew
rlabel metal3 s 27705 4903 27803 5001 4 vdd
port 2 nsew
rlabel metal3 s 32584 2513 32682 2611 4 vdd
port 2 nsew
rlabel metal3 s 32604 1563 32702 1661 4 vdd
port 2 nsew
rlabel metal3 s 27717 4065 27815 4163 4 vdd
port 2 nsew
rlabel metal3 s 30456 7426 30554 7524 4 gnd
port 3 nsew
rlabel metal3 s 31356 1563 31454 1661 4 vdd
port 2 nsew
rlabel metal3 s 31457 2181 31555 2279 4 gnd
port 3 nsew
rlabel metal3 s 27592 2513 27690 2611 4 vdd
port 2 nsew
rlabel metal3 s 30213 4065 30311 4163 4 vdd
port 2 nsew
rlabel metal3 s 26457 4903 26555 5001 4 vdd
port 2 nsew
rlabel metal3 s 28961 2181 29059 2279 4 gnd
port 3 nsew
rlabel metal3 s 27717 3743 27815 3841 4 gnd
port 3 nsew
rlabel metal3 s 30088 2513 30186 2611 4 vdd
port 2 nsew
rlabel metal3 s 28846 1979 28944 2077 4 gnd
port 3 nsew
rlabel metal3 s 27598 1979 27696 2077 4 gnd
port 3 nsew
rlabel metal3 s 28851 2950 28949 3048 4 gnd
port 3 nsew
rlabel metal3 s 27713 2181 27811 2279 4 gnd
port 3 nsew
rlabel metal3 s 26350 1979 26448 2077 4 gnd
port 3 nsew
rlabel metal3 s 30094 1979 30192 2077 4 gnd
port 3 nsew
rlabel metal3 s 30201 4903 30299 5001 4 vdd
port 2 nsew
rlabel metal3 s 31347 2950 31445 3048 4 gnd
port 3 nsew
rlabel metal3 s 27603 2950 27701 3048 4 gnd
port 3 nsew
rlabel metal3 s 31531 5677 31629 5775 4 gnd
port 3 nsew
rlabel metal3 s 29208 7426 29306 7524 4 gnd
port 3 nsew
rlabel metal3 s 32590 1979 32688 2077 4 gnd
port 3 nsew
rlabel metal3 s 27787 5677 27885 5775 4 gnd
port 3 nsew
rlabel metal3 s 31336 2513 31434 2611 4 vdd
port 2 nsew
rlabel metal3 s 32952 7426 33050 7524 4 gnd
port 3 nsew
rlabel metal3 s 32705 2181 32803 2279 4 gnd
port 3 nsew
rlabel metal3 s 31461 4065 31559 4163 4 vdd
port 2 nsew
rlabel metal3 s 31449 4903 31547 5001 4 vdd
port 2 nsew
rlabel metal3 s 32709 4065 32807 4163 4 vdd
port 2 nsew
rlabel metal3 s 30108 1563 30206 1661 4 vdd
port 2 nsew
rlabel metal3 s 26469 4065 26567 4163 4 vdd
port 2 nsew
rlabel metal3 s 32709 3743 32807 3841 4 gnd
port 3 nsew
rlabel metal3 s 31342 1979 31440 2077 4 gnd
port 3 nsew
rlabel metal3 s 29035 5677 29133 5775 4 gnd
port 3 nsew
rlabel metal3 s 28965 3743 29063 3841 4 gnd
port 3 nsew
rlabel metal3 s 30099 2950 30197 3048 4 gnd
port 3 nsew
rlabel metal3 s 32595 2950 32693 3048 4 gnd
port 3 nsew
rlabel metal3 s 28953 4903 29051 5001 4 vdd
port 2 nsew
rlabel metal3 s 26712 7426 26810 7524 4 gnd
port 3 nsew
rlabel metal3 s 26344 2513 26442 2611 4 vdd
port 2 nsew
rlabel metal3 s 26355 2950 26453 3048 4 gnd
port 3 nsew
rlabel metal3 s 28965 4065 29063 4163 4 vdd
port 2 nsew
rlabel metal3 s 26465 2181 26563 2279 4 gnd
port 3 nsew
rlabel metal3 s 30209 2181 30307 2279 4 gnd
port 3 nsew
rlabel metal3 s 28840 2513 28938 2611 4 vdd
port 2 nsew
rlabel metal3 s 26539 5677 26637 5775 4 gnd
port 3 nsew
rlabel metal3 s 26364 1563 26462 1661 4 vdd
port 2 nsew
rlabel metal3 s 30283 5677 30381 5775 4 gnd
port 3 nsew
rlabel metal3 s 32697 4903 32795 5001 4 vdd
port 2 nsew
rlabel metal3 s 27960 7426 28058 7524 4 gnd
port 3 nsew
rlabel metal3 s 31461 3743 31559 3841 4 gnd
port 3 nsew
rlabel metal3 s 28860 1563 28958 1661 4 vdd
port 2 nsew
rlabel metal3 s 31704 7426 31802 7524 4 gnd
port 3 nsew
rlabel metal3 s 30213 3743 30311 3841 4 gnd
port 3 nsew
rlabel metal3 s 32779 5677 32877 5775 4 gnd
port 3 nsew
rlabel metal3 s 60702 32233 60800 32331 4 vdd
port 2 nsew
rlabel metal3 s 60270 29505 60368 29603 4 vdd
port 2 nsew
rlabel metal3 s 60270 29863 60368 29961 4 vdd
port 2 nsew
rlabel metal3 s 60702 29863 60800 29961 4 vdd
port 2 nsew
rlabel metal3 s 61127 31501 61225 31599 4 gnd
port 3 nsew
rlabel metal3 s 60702 29505 60800 29603 4 vdd
port 2 nsew
rlabel metal3 s 59888 30272 59986 30370 4 gnd
port 3 nsew
rlabel metal3 s 59492 29877 59590 29975 4 vdd
port 2 nsew
rlabel metal3 s 60270 31875 60368 31973 4 vdd
port 2 nsew
rlabel metal3 s 60702 31875 60800 31973 4 vdd
port 2 nsew
rlabel metal3 s 60702 30653 60800 30751 4 vdd
port 2 nsew
rlabel metal3 s 59492 30667 59590 30765 4 vdd
port 2 nsew
rlabel metal3 s 60270 31085 60368 31183 4 vdd
port 2 nsew
rlabel metal3 s 61127 33081 61225 33179 4 gnd
port 3 nsew
rlabel metal3 s 59888 29877 59986 29975 4 gnd
port 3 nsew
rlabel metal3 s 59888 33432 59986 33530 4 gnd
port 3 nsew
rlabel metal3 s 61127 29505 61225 29603 4 gnd
port 3 nsew
rlabel metal3 s 59492 33432 59590 33530 4 vdd
port 2 nsew
rlabel metal3 s 59492 31457 59590 31555 4 vdd
port 2 nsew
rlabel metal3 s 60270 30653 60368 30751 4 vdd
port 2 nsew
rlabel metal3 s 60270 31443 60368 31541 4 vdd
port 2 nsew
rlabel metal3 s 60270 33023 60368 33121 4 vdd
port 2 nsew
rlabel metal3 s 60702 31085 60800 31183 4 vdd
port 2 nsew
rlabel metal3 s 59492 31062 59590 31160 4 vdd
port 2 nsew
rlabel metal3 s 59888 31852 59986 31950 4 gnd
port 3 nsew
rlabel metal3 s 60270 33455 60368 33553 4 vdd
port 2 nsew
rlabel metal3 s 60702 33455 60800 33553 4 vdd
port 2 nsew
rlabel metal3 s 59888 29482 59986 29580 4 gnd
port 3 nsew
rlabel metal3 s 61127 30711 61225 30809 4 gnd
port 3 nsew
rlabel metal3 s 60702 30295 60800 30393 4 vdd
port 2 nsew
rlabel metal3 s 60702 32665 60800 32763 4 vdd
port 2 nsew
rlabel metal3 s 60270 32233 60368 32331 4 vdd
port 2 nsew
rlabel metal3 s 59888 33037 59986 33135 4 gnd
port 3 nsew
rlabel metal3 s 59888 31062 59986 31160 4 gnd
port 3 nsew
rlabel metal3 s 59492 30272 59590 30370 4 vdd
port 2 nsew
rlabel metal3 s 60270 32665 60368 32763 4 vdd
port 2 nsew
rlabel metal3 s 59492 29482 59590 29580 4 vdd
port 2 nsew
rlabel metal3 s 61127 32291 61225 32389 4 gnd
port 3 nsew
rlabel metal3 s 59888 31457 59986 31555 4 gnd
port 3 nsew
rlabel metal3 s 59492 32247 59590 32345 4 vdd
port 2 nsew
rlabel metal3 s 59492 33037 59590 33135 4 vdd
port 2 nsew
rlabel metal3 s 60702 33023 60800 33121 4 vdd
port 2 nsew
rlabel metal3 s 61127 29921 61225 30019 4 gnd
port 3 nsew
rlabel metal3 s 61127 31085 61225 31183 4 gnd
port 3 nsew
rlabel metal3 s 61127 30295 61225 30393 4 gnd
port 3 nsew
rlabel metal3 s 60702 31443 60800 31541 4 vdd
port 2 nsew
rlabel metal3 s 60270 30295 60368 30393 4 vdd
port 2 nsew
rlabel metal3 s 59492 31852 59590 31950 4 vdd
port 2 nsew
rlabel metal3 s 61127 31875 61225 31973 4 gnd
port 3 nsew
rlabel metal3 s 59888 32642 59986 32740 4 gnd
port 3 nsew
rlabel metal3 s 61127 33455 61225 33553 4 gnd
port 3 nsew
rlabel metal3 s 59492 32642 59590 32740 4 vdd
port 2 nsew
rlabel metal3 s 59888 30667 59986 30765 4 gnd
port 3 nsew
rlabel metal3 s 61127 32665 61225 32763 4 gnd
port 3 nsew
rlabel metal3 s 59888 32247 59986 32345 4 gnd
port 3 nsew
rlabel metal3 s 59888 27507 59986 27605 4 gnd
port 3 nsew
rlabel metal3 s 61127 27925 61225 28023 4 gnd
port 3 nsew
rlabel metal3 s 60702 27925 60800 28023 4 vdd
port 2 nsew
rlabel metal3 s 61127 28341 61225 28439 4 gnd
port 3 nsew
rlabel metal3 s 59492 26717 59590 26815 4 vdd
port 2 nsew
rlabel metal3 s 61127 25555 61225 25653 4 gnd
port 3 nsew
rlabel metal3 s 61127 27135 61225 27233 4 gnd
port 3 nsew
rlabel metal3 s 60702 25555 60800 25653 4 vdd
port 2 nsew
rlabel metal3 s 59492 29087 59590 29185 4 vdd
port 2 nsew
rlabel metal3 s 59492 27902 59590 28000 4 vdd
port 2 nsew
rlabel metal3 s 60270 29073 60368 29171 4 vdd
port 2 nsew
rlabel metal3 s 60702 26703 60800 26801 4 vdd
port 2 nsew
rlabel metal3 s 60270 28283 60368 28381 4 vdd
port 2 nsew
rlabel metal3 s 59492 25927 59590 26025 4 vdd
port 2 nsew
rlabel metal3 s 60702 29073 60800 29171 4 vdd
port 2 nsew
rlabel metal3 s 60702 26345 60800 26443 4 vdd
port 2 nsew
rlabel metal3 s 59492 25532 59590 25630 4 vdd
port 2 nsew
rlabel metal3 s 61127 27551 61225 27649 4 gnd
port 3 nsew
rlabel metal3 s 59888 25927 59986 26025 4 gnd
port 3 nsew
rlabel metal3 s 60270 27135 60368 27233 4 vdd
port 2 nsew
rlabel metal3 s 61127 25181 61225 25279 4 gnd
port 3 nsew
rlabel metal3 s 59888 28692 59986 28790 4 gnd
port 3 nsew
rlabel metal3 s 61127 28715 61225 28813 4 gnd
port 3 nsew
rlabel metal3 s 59888 28297 59986 28395 4 gnd
port 3 nsew
rlabel metal3 s 59492 27112 59590 27210 4 vdd
port 2 nsew
rlabel metal3 s 59888 29087 59986 29185 4 gnd
port 3 nsew
rlabel metal3 s 61127 29131 61225 29229 4 gnd
port 3 nsew
rlabel metal3 s 59492 26322 59590 26420 4 vdd
port 2 nsew
rlabel metal3 s 59492 28692 59590 28790 4 vdd
port 2 nsew
rlabel metal3 s 59888 25532 59986 25630 4 gnd
port 3 nsew
rlabel metal3 s 60702 28715 60800 28813 4 vdd
port 2 nsew
rlabel metal3 s 59888 27112 59986 27210 4 gnd
port 3 nsew
rlabel metal3 s 60270 25913 60368 26011 4 vdd
port 2 nsew
rlabel metal3 s 60702 27135 60800 27233 4 vdd
port 2 nsew
rlabel metal3 s 59492 28297 59590 28395 4 vdd
port 2 nsew
rlabel metal3 s 60270 26345 60368 26443 4 vdd
port 2 nsew
rlabel metal3 s 59888 27902 59986 28000 4 gnd
port 3 nsew
rlabel metal3 s 60702 25913 60800 26011 4 vdd
port 2 nsew
rlabel metal3 s 59888 26322 59986 26420 4 gnd
port 3 nsew
rlabel metal3 s 59492 27507 59590 27605 4 vdd
port 2 nsew
rlabel metal3 s 59888 26717 59986 26815 4 gnd
port 3 nsew
rlabel metal3 s 60270 26703 60368 26801 4 vdd
port 2 nsew
rlabel metal3 s 60270 25555 60368 25653 4 vdd
port 2 nsew
rlabel metal3 s 61127 26345 61225 26443 4 gnd
port 3 nsew
rlabel metal3 s 61127 26761 61225 26859 4 gnd
port 3 nsew
rlabel metal3 s 60702 27493 60800 27591 4 vdd
port 2 nsew
rlabel metal3 s 60270 27925 60368 28023 4 vdd
port 2 nsew
rlabel metal3 s 60270 27493 60368 27591 4 vdd
port 2 nsew
rlabel metal3 s 61127 25971 61225 26069 4 gnd
port 3 nsew
rlabel metal3 s 60270 28715 60368 28813 4 vdd
port 2 nsew
rlabel metal3 s 60702 28283 60800 28381 4 vdd
port 2 nsew
rlabel metal3 s 54552 26717 54650 26815 4 gnd
port 3 nsew
rlabel metal3 s 54552 25927 54650 26025 4 gnd
port 3 nsew
rlabel metal3 s 54552 29324 54650 29422 4 gnd
port 3 nsew
rlabel metal3 s 54552 27744 54650 27842 4 gnd
port 3 nsew
rlabel metal3 s 54552 29877 54650 29975 4 gnd
port 3 nsew
rlabel metal3 s 54552 30114 54650 30212 4 gnd
port 3 nsew
rlabel metal3 s 54552 28534 54650 28632 4 gnd
port 3 nsew
rlabel metal3 s 54552 25374 54650 25472 4 gnd
port 3 nsew
rlabel metal3 s 54552 27270 54650 27368 4 gnd
port 3 nsew
rlabel metal3 s 54552 32010 54650 32108 4 gnd
port 3 nsew
rlabel metal3 s 54552 26164 54650 26262 4 gnd
port 3 nsew
rlabel metal3 s 54552 33037 54650 33135 4 gnd
port 3 nsew
rlabel metal3 s 54552 30430 54650 30528 4 gnd
port 3 nsew
rlabel metal3 s 54552 31220 54650 31318 4 gnd
port 3 nsew
rlabel metal3 s 54552 33274 54650 33372 4 gnd
port 3 nsew
rlabel metal3 s 54552 28297 54650 28395 4 gnd
port 3 nsew
rlabel metal3 s 54552 27507 54650 27605 4 gnd
port 3 nsew
rlabel metal3 s 54552 28060 54650 28158 4 gnd
port 3 nsew
rlabel metal3 s 54552 28850 54650 28948 4 gnd
port 3 nsew
rlabel metal3 s 54552 31694 54650 31792 4 gnd
port 3 nsew
rlabel metal3 s 54552 26954 54650 27052 4 gnd
port 3 nsew
rlabel metal3 s 54552 30667 54650 30765 4 gnd
port 3 nsew
rlabel metal3 s 54552 29087 54650 29185 4 gnd
port 3 nsew
rlabel metal3 s 54552 32800 54650 32898 4 gnd
port 3 nsew
rlabel metal3 s 54552 31457 54650 31555 4 gnd
port 3 nsew
rlabel metal3 s 54552 32484 54650 32582 4 gnd
port 3 nsew
rlabel metal3 s 54552 29640 54650 29738 4 gnd
port 3 nsew
rlabel metal3 s 54552 26480 54650 26578 4 gnd
port 3 nsew
rlabel metal3 s 54552 30904 54650 31002 4 gnd
port 3 nsew
rlabel metal3 s 54552 32247 54650 32345 4 gnd
port 3 nsew
rlabel metal3 s 54552 25690 54650 25788 4 gnd
port 3 nsew
rlabel metal3 s 54552 21187 54650 21285 4 gnd
port 3 nsew
rlabel metal3 s 54552 21424 54650 21522 4 gnd
port 3 nsew
rlabel metal3 s 54552 18027 54650 18125 4 gnd
port 3 nsew
rlabel metal3 s 54552 17000 54650 17098 4 gnd
port 3 nsew
rlabel metal3 s 54552 19370 54650 19468 4 gnd
port 3 nsew
rlabel metal3 s 54552 18817 54650 18915 4 gnd
port 3 nsew
rlabel metal3 s 54552 25137 54650 25235 4 gnd
port 3 nsew
rlabel metal3 s 54552 21740 54650 21838 4 gnd
port 3 nsew
rlabel metal3 s 54552 20634 54650 20732 4 gnd
port 3 nsew
rlabel metal3 s 54552 17790 54650 17888 4 gnd
port 3 nsew
rlabel metal3 s 54552 23557 54650 23655 4 gnd
port 3 nsew
rlabel metal3 s 54552 19054 54650 19152 4 gnd
port 3 nsew
rlabel metal3 s 54552 24347 54650 24445 4 gnd
port 3 nsew
rlabel metal3 s 54552 23794 54650 23892 4 gnd
port 3 nsew
rlabel metal3 s 54552 24900 54650 24998 4 gnd
port 3 nsew
rlabel metal3 s 54552 19607 54650 19705 4 gnd
port 3 nsew
rlabel metal3 s 54552 21977 54650 22075 4 gnd
port 3 nsew
rlabel metal3 s 54552 19844 54650 19942 4 gnd
port 3 nsew
rlabel metal3 s 54552 22530 54650 22628 4 gnd
port 3 nsew
rlabel metal3 s 54552 22767 54650 22865 4 gnd
port 3 nsew
rlabel metal3 s 54552 18264 54650 18362 4 gnd
port 3 nsew
rlabel metal3 s 54552 24110 54650 24208 4 gnd
port 3 nsew
rlabel metal3 s 54552 23320 54650 23418 4 gnd
port 3 nsew
rlabel metal3 s 54552 20950 54650 21048 4 gnd
port 3 nsew
rlabel metal3 s 54552 17237 54650 17335 4 gnd
port 3 nsew
rlabel metal3 s 54552 23004 54650 23102 4 gnd
port 3 nsew
rlabel metal3 s 54552 18580 54650 18678 4 gnd
port 3 nsew
rlabel metal3 s 54552 20397 54650 20495 4 gnd
port 3 nsew
rlabel metal3 s 54552 22214 54650 22312 4 gnd
port 3 nsew
rlabel metal3 s 54552 20160 54650 20258 4 gnd
port 3 nsew
rlabel metal3 s 54552 17474 54650 17572 4 gnd
port 3 nsew
rlabel metal3 s 54552 24584 54650 24682 4 gnd
port 3 nsew
rlabel metal3 s 60270 22753 60368 22851 4 vdd
port 2 nsew
rlabel metal3 s 61127 21605 61225 21703 4 gnd
port 3 nsew
rlabel metal3 s 59492 24742 59590 24840 4 vdd
port 2 nsew
rlabel metal3 s 60270 21605 60368 21703 4 vdd
port 2 nsew
rlabel metal3 s 60702 23975 60800 24073 4 vdd
port 2 nsew
rlabel metal3 s 59888 22372 59986 22470 4 gnd
port 3 nsew
rlabel metal3 s 61127 21231 61225 21329 4 gnd
port 3 nsew
rlabel metal3 s 60270 23185 60368 23283 4 vdd
port 2 nsew
rlabel metal3 s 60270 25123 60368 25221 4 vdd
port 2 nsew
rlabel metal3 s 59492 21187 59590 21285 4 vdd
port 2 nsew
rlabel metal3 s 60702 21963 60800 22061 4 vdd
port 2 nsew
rlabel metal3 s 61127 24765 61225 24863 4 gnd
port 3 nsew
rlabel metal3 s 60270 21963 60368 22061 4 vdd
port 2 nsew
rlabel metal3 s 59492 21977 59590 22075 4 vdd
port 2 nsew
rlabel metal3 s 60702 24765 60800 24863 4 vdd
port 2 nsew
rlabel metal3 s 59888 24347 59986 24445 4 gnd
port 3 nsew
rlabel metal3 s 60270 22395 60368 22493 4 vdd
port 2 nsew
rlabel metal3 s 59888 23952 59986 24050 4 gnd
port 3 nsew
rlabel metal3 s 60270 21173 60368 21271 4 vdd
port 2 nsew
rlabel metal3 s 59492 23952 59590 24050 4 vdd
port 2 nsew
rlabel metal3 s 60702 22395 60800 22493 4 vdd
port 2 nsew
rlabel metal3 s 59888 23162 59986 23260 4 gnd
port 3 nsew
rlabel metal3 s 60270 23975 60368 24073 4 vdd
port 2 nsew
rlabel metal3 s 61127 22021 61225 22119 4 gnd
port 3 nsew
rlabel metal3 s 60702 21173 60800 21271 4 vdd
port 2 nsew
rlabel metal3 s 60702 23543 60800 23641 4 vdd
port 2 nsew
rlabel metal3 s 59888 23557 59986 23655 4 gnd
port 3 nsew
rlabel metal3 s 60270 24333 60368 24431 4 vdd
port 2 nsew
rlabel metal3 s 59492 22372 59590 22470 4 vdd
port 2 nsew
rlabel metal3 s 59492 25137 59590 25235 4 vdd
port 2 nsew
rlabel metal3 s 59888 24742 59986 24840 4 gnd
port 3 nsew
rlabel metal3 s 60702 22753 60800 22851 4 vdd
port 2 nsew
rlabel metal3 s 59888 21187 59986 21285 4 gnd
port 3 nsew
rlabel metal3 s 59492 23557 59590 23655 4 vdd
port 2 nsew
rlabel metal3 s 61127 24391 61225 24489 4 gnd
port 3 nsew
rlabel metal3 s 61127 23601 61225 23699 4 gnd
port 3 nsew
rlabel metal3 s 60702 25123 60800 25221 4 vdd
port 2 nsew
rlabel metal3 s 60270 24765 60368 24863 4 vdd
port 2 nsew
rlabel metal3 s 59888 21977 59986 22075 4 gnd
port 3 nsew
rlabel metal3 s 59492 24347 59590 24445 4 vdd
port 2 nsew
rlabel metal3 s 61127 23185 61225 23283 4 gnd
port 3 nsew
rlabel metal3 s 59492 22767 59590 22865 4 vdd
port 2 nsew
rlabel metal3 s 60270 23543 60368 23641 4 vdd
port 2 nsew
rlabel metal3 s 59492 23162 59590 23260 4 vdd
port 2 nsew
rlabel metal3 s 61127 22811 61225 22909 4 gnd
port 3 nsew
rlabel metal3 s 59888 21582 59986 21680 4 gnd
port 3 nsew
rlabel metal3 s 60702 23185 60800 23283 4 vdd
port 2 nsew
rlabel metal3 s 60702 21605 60800 21703 4 vdd
port 2 nsew
rlabel metal3 s 59888 25137 59986 25235 4 gnd
port 3 nsew
rlabel metal3 s 61127 22395 61225 22493 4 gnd
port 3 nsew
rlabel metal3 s 59492 21582 59590 21680 4 vdd
port 2 nsew
rlabel metal3 s 61127 23975 61225 24073 4 gnd
port 3 nsew
rlabel metal3 s 60702 24333 60800 24431 4 vdd
port 2 nsew
rlabel metal3 s 59888 22767 59986 22865 4 gnd
port 3 nsew
rlabel metal3 s 60270 19235 60368 19333 4 vdd
port 2 nsew
rlabel metal3 s 60702 17223 60800 17321 4 vdd
port 2 nsew
rlabel metal3 s 60270 19593 60368 19691 4 vdd
port 2 nsew
rlabel metal3 s 60702 20815 60800 20913 4 vdd
port 2 nsew
rlabel metal3 s 61127 20815 61225 20913 4 gnd
port 3 nsew
rlabel metal3 s 60702 19593 60800 19691 4 vdd
port 2 nsew
rlabel metal3 s 60702 18445 60800 18543 4 vdd
port 2 nsew
rlabel metal3 s 61127 17655 61225 17753 4 gnd
port 3 nsew
rlabel metal3 s 59492 18422 59590 18520 4 vdd
port 2 nsew
rlabel metal3 s 60270 20815 60368 20913 4 vdd
port 2 nsew
rlabel metal3 s 59492 19212 59590 19310 4 vdd
port 2 nsew
rlabel metal3 s 59888 16842 59986 16940 4 gnd
port 3 nsew
rlabel metal3 s 59888 17632 59986 17730 4 gnd
port 3 nsew
rlabel metal3 s 60702 16865 60800 16963 4 vdd
port 2 nsew
rlabel metal3 s 59888 19607 59986 19705 4 gnd
port 3 nsew
rlabel metal3 s 60270 16865 60368 16963 4 vdd
port 2 nsew
rlabel metal3 s 59492 20792 59590 20890 4 vdd
port 2 nsew
rlabel metal3 s 59492 17632 59590 17730 4 vdd
port 2 nsew
rlabel metal3 s 60270 18013 60368 18111 4 vdd
port 2 nsew
rlabel metal3 s 59888 18422 59986 18520 4 gnd
port 3 nsew
rlabel metal3 s 59492 18027 59590 18125 4 vdd
port 2 nsew
rlabel metal3 s 59888 20397 59986 20495 4 gnd
port 3 nsew
rlabel metal3 s 61127 20441 61225 20539 4 gnd
port 3 nsew
rlabel metal3 s 61127 19651 61225 19749 4 gnd
port 3 nsew
rlabel metal3 s 60702 19235 60800 19333 4 vdd
port 2 nsew
rlabel metal3 s 59492 20397 59590 20495 4 vdd
port 2 nsew
rlabel metal3 s 59888 18817 59986 18915 4 gnd
port 3 nsew
rlabel metal3 s 61127 16865 61225 16963 4 gnd
port 3 nsew
rlabel metal3 s 59888 20002 59986 20100 4 gnd
port 3 nsew
rlabel metal3 s 59888 17237 59986 17335 4 gnd
port 3 nsew
rlabel metal3 s 60702 20025 60800 20123 4 vdd
port 2 nsew
rlabel metal3 s 61127 17281 61225 17379 4 gnd
port 3 nsew
rlabel metal3 s 60270 18445 60368 18543 4 vdd
port 2 nsew
rlabel metal3 s 61127 18445 61225 18543 4 gnd
port 3 nsew
rlabel metal3 s 61127 20025 61225 20123 4 gnd
port 3 nsew
rlabel metal3 s 60270 20383 60368 20481 4 vdd
port 2 nsew
rlabel metal3 s 60270 18803 60368 18901 4 vdd
port 2 nsew
rlabel metal3 s 59492 17237 59590 17335 4 vdd
port 2 nsew
rlabel metal3 s 61127 19235 61225 19333 4 gnd
port 3 nsew
rlabel metal3 s 61127 18071 61225 18169 4 gnd
port 3 nsew
rlabel metal3 s 60702 20383 60800 20481 4 vdd
port 2 nsew
rlabel metal3 s 60702 18803 60800 18901 4 vdd
port 2 nsew
rlabel metal3 s 60270 17655 60368 17753 4 vdd
port 2 nsew
rlabel metal3 s 59492 20002 59590 20100 4 vdd
port 2 nsew
rlabel metal3 s 59888 18027 59986 18125 4 gnd
port 3 nsew
rlabel metal3 s 59492 19607 59590 19705 4 vdd
port 2 nsew
rlabel metal3 s 60702 18013 60800 18111 4 vdd
port 2 nsew
rlabel metal3 s 61127 18861 61225 18959 4 gnd
port 3 nsew
rlabel metal3 s 59492 18817 59590 18915 4 vdd
port 2 nsew
rlabel metal3 s 60270 20025 60368 20123 4 vdd
port 2 nsew
rlabel metal3 s 60702 17655 60800 17753 4 vdd
port 2 nsew
rlabel metal3 s 59888 19212 59986 19310 4 gnd
port 3 nsew
rlabel metal3 s 59492 16842 59590 16940 4 vdd
port 2 nsew
rlabel metal3 s 60270 17223 60368 17321 4 vdd
port 2 nsew
rlabel metal3 s 59888 20792 59986 20890 4 gnd
port 3 nsew
rlabel metal3 s 64541 16865 64639 16963 4 gnd
port 3 nsew
rlabel metal3 s 63684 17655 63782 17753 4 vdd
port 2 nsew
rlabel metal3 s 62906 17632 63004 17730 4 vdd
port 2 nsew
rlabel metal3 s 63302 16842 63400 16940 4 gnd
port 3 nsew
rlabel metal3 s 64116 17655 64214 17753 4 vdd
port 2 nsew
rlabel metal3 s 63684 16865 63782 16963 4 vdd
port 2 nsew
rlabel metal3 s 63302 17632 63400 17730 4 gnd
port 3 nsew
rlabel metal3 s 64116 16865 64214 16963 4 vdd
port 2 nsew
rlabel metal3 s 64541 17655 64639 17753 4 gnd
port 3 nsew
rlabel metal3 s 62906 16842 63004 16940 4 vdd
port 2 nsew
rlabel metal3 s 48240 9566 48338 9664 4 vdd
port 2 nsew
rlabel metal3 s 45001 8975 45099 9073 4 vdd
port 2 nsew
rlabel metal3 s 49607 8975 49705 9073 4 vdd
port 2 nsew
rlabel metal3 s 43872 9566 43970 9664 4 vdd
port 2 nsew
rlabel metal3 s 48864 9566 48962 9664 4 vdd
port 2 nsew
rlabel metal3 s 46249 8975 46347 9073 4 vdd
port 2 nsew
rlabel metal3 s 42000 9566 42098 9664 4 vdd
port 2 nsew
rlabel metal3 s 43248 9566 43346 9664 4 vdd
port 2 nsew
rlabel metal3 s 42119 8975 42217 9073 4 vdd
port 2 nsew
rlabel metal3 s 42505 8975 42603 9073 4 vdd
port 2 nsew
rlabel metal3 s 48359 8975 48457 9073 4 vdd
port 2 nsew
rlabel metal3 s 47497 8975 47595 9073 4 vdd
port 2 nsew
rlabel metal3 s 43753 8975 43851 9073 4 vdd
port 2 nsew
rlabel metal3 s 47616 9566 47714 9664 4 vdd
port 2 nsew
rlabel metal3 s 49488 9566 49586 9664 4 vdd
port 2 nsew
rlabel metal3 s 46368 9566 46466 9664 4 vdd
port 2 nsew
rlabel metal3 s 43367 8975 43465 9073 4 vdd
port 2 nsew
rlabel metal3 s 46992 9566 47090 9664 4 vdd
port 2 nsew
rlabel metal3 s 47111 8975 47209 9073 4 vdd
port 2 nsew
rlabel metal3 s 44615 8975 44713 9073 4 vdd
port 2 nsew
rlabel metal3 s 44496 9566 44594 9664 4 vdd
port 2 nsew
rlabel metal3 s 48745 8975 48843 9073 4 vdd
port 2 nsew
rlabel metal3 s 42624 9566 42722 9664 4 vdd
port 2 nsew
rlabel metal3 s 45863 8975 45961 9073 4 vdd
port 2 nsew
rlabel metal3 s 45120 9566 45218 9664 4 vdd
port 2 nsew
rlabel metal3 s 45744 9566 45842 9664 4 vdd
port 2 nsew
rlabel metal3 s 40128 9566 40226 9664 4 vdd
port 2 nsew
rlabel metal3 s 41376 9566 41474 9664 4 vdd
port 2 nsew
rlabel metal3 s 39623 8975 39721 9073 4 vdd
port 2 nsew
rlabel metal3 s 37632 9566 37730 9664 4 vdd
port 2 nsew
rlabel metal3 s 38256 9566 38354 9664 4 vdd
port 2 nsew
rlabel metal3 s 37127 8975 37225 9073 4 vdd
port 2 nsew
rlabel metal3 s 37513 8975 37611 9073 4 vdd
port 2 nsew
rlabel metal3 s 38375 8975 38473 9073 4 vdd
port 2 nsew
rlabel metal3 s 34631 8975 34729 9073 4 vdd
port 2 nsew
rlabel metal3 s 41257 8975 41355 9073 4 vdd
port 2 nsew
rlabel metal3 s 33769 8975 33867 9073 4 vdd
port 2 nsew
rlabel metal3 s 35136 9566 35234 9664 4 vdd
port 2 nsew
rlabel metal3 s 40752 9566 40850 9664 4 vdd
port 2 nsew
rlabel metal3 s 36265 8975 36363 9073 4 vdd
port 2 nsew
rlabel metal3 s 40871 8975 40969 9073 4 vdd
port 2 nsew
rlabel metal3 s 33888 9566 33986 9664 4 vdd
port 2 nsew
rlabel metal3 s 35879 8975 35977 9073 4 vdd
port 2 nsew
rlabel metal3 s 37008 9566 37106 9664 4 vdd
port 2 nsew
rlabel metal3 s 35760 9566 35858 9664 4 vdd
port 2 nsew
rlabel metal3 s 34512 9566 34610 9664 4 vdd
port 2 nsew
rlabel metal3 s 38880 9566 38978 9664 4 vdd
port 2 nsew
rlabel metal3 s 36384 9566 36482 9664 4 vdd
port 2 nsew
rlabel metal3 s 35017 8975 35115 9073 4 vdd
port 2 nsew
rlabel metal3 s 40009 8975 40107 9073 4 vdd
port 2 nsew
rlabel metal3 s 39504 9566 39602 9664 4 vdd
port 2 nsew
rlabel metal3 s 38761 8975 38859 9073 4 vdd
port 2 nsew
rlabel metal3 s 40440 7426 40538 7524 4 gnd
port 3 nsew
rlabel metal3 s 41515 5677 41613 5775 4 gnd
port 3 nsew
rlabel metal3 s 38830 1979 38928 2077 4 gnd
port 3 nsew
rlabel metal3 s 37582 1979 37680 2077 4 gnd
port 3 nsew
rlabel metal3 s 35086 1979 35184 2077 4 gnd
port 3 nsew
rlabel metal3 s 41326 1979 41424 2077 4 gnd
port 3 nsew
rlabel metal3 s 35275 5677 35373 5775 4 gnd
port 3 nsew
rlabel metal3 s 33957 4065 34055 4163 4 vdd
port 2 nsew
rlabel metal3 s 36339 2950 36437 3048 4 gnd
port 3 nsew
rlabel metal3 s 36441 4903 36539 5001 4 vdd
port 2 nsew
rlabel metal3 s 36696 7426 36794 7524 4 gnd
port 3 nsew
rlabel metal3 s 35448 7426 35546 7524 4 gnd
port 3 nsew
rlabel metal3 s 40197 3743 40295 3841 4 gnd
port 3 nsew
rlabel metal3 s 38835 2950 38933 3048 4 gnd
port 3 nsew
rlabel metal3 s 38945 2181 39043 2279 4 gnd
port 3 nsew
rlabel metal3 s 40185 4903 40283 5001 4 vdd
port 2 nsew
rlabel metal3 s 34027 5677 34125 5775 4 gnd
port 3 nsew
rlabel metal3 s 40193 2181 40291 2279 4 gnd
port 3 nsew
rlabel metal3 s 38937 4903 39035 5001 4 vdd
port 2 nsew
rlabel metal3 s 35100 1563 35198 1661 4 vdd
port 2 nsew
rlabel metal3 s 40267 5677 40365 5775 4 gnd
port 3 nsew
rlabel metal3 s 40083 2950 40181 3048 4 gnd
port 3 nsew
rlabel metal3 s 34200 7426 34298 7524 4 gnd
port 3 nsew
rlabel metal3 s 36328 2513 36426 2611 4 vdd
port 2 nsew
rlabel metal3 s 37771 5677 37869 5775 4 gnd
port 3 nsew
rlabel metal3 s 38949 4065 39047 4163 4 vdd
port 2 nsew
rlabel metal3 s 36453 3743 36551 3841 4 gnd
port 3 nsew
rlabel metal3 s 33843 2950 33941 3048 4 gnd
port 3 nsew
rlabel metal3 s 35205 3743 35303 3841 4 gnd
port 3 nsew
rlabel metal3 s 33945 4903 34043 5001 4 vdd
port 2 nsew
rlabel metal3 s 39192 7426 39290 7524 4 gnd
port 3 nsew
rlabel metal3 s 35091 2950 35189 3048 4 gnd
port 3 nsew
rlabel metal3 s 41445 4065 41543 4163 4 vdd
port 2 nsew
rlabel metal3 s 35193 4903 35291 5001 4 vdd
port 2 nsew
rlabel metal3 s 40092 1563 40190 1661 4 vdd
port 2 nsew
rlabel metal3 s 41433 4903 41531 5001 4 vdd
port 2 nsew
rlabel metal3 s 40197 4065 40295 4163 4 vdd
port 2 nsew
rlabel metal3 s 37944 7426 38042 7524 4 gnd
port 3 nsew
rlabel metal3 s 40078 1979 40176 2077 4 gnd
port 3 nsew
rlabel metal3 s 37596 1563 37694 1661 4 vdd
port 2 nsew
rlabel metal3 s 35080 2513 35178 2611 4 vdd
port 2 nsew
rlabel metal3 s 36334 1979 36432 2077 4 gnd
port 3 nsew
rlabel metal3 s 41331 2950 41429 3048 4 gnd
port 3 nsew
rlabel metal3 s 36453 4065 36551 4163 4 vdd
port 2 nsew
rlabel metal3 s 39019 5677 39117 5775 4 gnd
port 3 nsew
rlabel metal3 s 40072 2513 40170 2611 4 vdd
port 2 nsew
rlabel metal3 s 36348 1563 36446 1661 4 vdd
port 2 nsew
rlabel metal3 s 38844 1563 38942 1661 4 vdd
port 2 nsew
rlabel metal3 s 37697 2181 37795 2279 4 gnd
port 3 nsew
rlabel metal3 s 41445 3743 41543 3841 4 gnd
port 3 nsew
rlabel metal3 s 37701 3743 37799 3841 4 gnd
port 3 nsew
rlabel metal3 s 38824 2513 38922 2611 4 vdd
port 2 nsew
rlabel metal3 s 41340 1563 41438 1661 4 vdd
port 2 nsew
rlabel metal3 s 36523 5677 36621 5775 4 gnd
port 3 nsew
rlabel metal3 s 41320 2513 41418 2611 4 vdd
port 2 nsew
rlabel metal3 s 33852 1563 33950 1661 4 vdd
port 2 nsew
rlabel metal3 s 38949 3743 39047 3841 4 gnd
port 3 nsew
rlabel metal3 s 36449 2181 36547 2279 4 gnd
port 3 nsew
rlabel metal3 s 33838 1979 33936 2077 4 gnd
port 3 nsew
rlabel metal3 s 33953 2181 34051 2279 4 gnd
port 3 nsew
rlabel metal3 s 37689 4903 37787 5001 4 vdd
port 2 nsew
rlabel metal3 s 37701 4065 37799 4163 4 vdd
port 2 nsew
rlabel metal3 s 41441 2181 41539 2279 4 gnd
port 3 nsew
rlabel metal3 s 33957 3743 34055 3841 4 gnd
port 3 nsew
rlabel metal3 s 35205 4065 35303 4163 4 vdd
port 2 nsew
rlabel metal3 s 37576 2513 37674 2611 4 vdd
port 2 nsew
rlabel metal3 s 33832 2513 33930 2611 4 vdd
port 2 nsew
rlabel metal3 s 35201 2181 35299 2279 4 gnd
port 3 nsew
rlabel metal3 s 37587 2950 37685 3048 4 gnd
port 3 nsew
rlabel metal3 s 48814 1979 48912 2077 4 gnd
port 3 nsew
rlabel metal3 s 47673 4903 47771 5001 4 vdd
port 2 nsew
rlabel metal3 s 47685 3743 47783 3841 4 gnd
port 3 nsew
rlabel metal3 s 43816 2513 43914 2611 4 vdd
port 2 nsew
rlabel metal3 s 47928 7426 48026 7524 4 gnd
port 3 nsew
rlabel metal3 s 45177 4903 45275 5001 4 vdd
port 2 nsew
rlabel metal3 s 45185 2181 45283 2279 4 gnd
port 3 nsew
rlabel metal3 s 47685 4065 47783 4163 4 vdd
port 2 nsew
rlabel metal3 s 46507 5677 46605 5775 4 gnd
port 3 nsew
rlabel metal3 s 45189 3743 45287 3841 4 gnd
port 3 nsew
rlabel metal3 s 44011 5677 44109 5775 4 gnd
port 3 nsew
rlabel metal3 s 47580 1563 47678 1661 4 vdd
port 2 nsew
rlabel metal3 s 48819 2950 48917 3048 4 gnd
port 3 nsew
rlabel metal3 s 45189 4065 45287 4163 4 vdd
port 2 nsew
rlabel metal3 s 45259 5677 45357 5775 4 gnd
port 3 nsew
rlabel metal3 s 45075 2950 45173 3048 4 gnd
port 3 nsew
rlabel metal3 s 48929 2181 49027 2279 4 gnd
port 3 nsew
rlabel metal3 s 43827 2950 43925 3048 4 gnd
port 3 nsew
rlabel metal3 s 48828 1563 48926 1661 4 vdd
port 2 nsew
rlabel metal3 s 42693 4065 42791 4163 4 vdd
port 2 nsew
rlabel metal3 s 43937 2181 44035 2279 4 gnd
port 3 nsew
rlabel metal3 s 46318 1979 46416 2077 4 gnd
port 3 nsew
rlabel metal3 s 42681 4903 42779 5001 4 vdd
port 2 nsew
rlabel metal3 s 47566 1979 47664 2077 4 gnd
port 3 nsew
rlabel metal3 s 48808 2513 48906 2611 4 vdd
port 2 nsew
rlabel metal3 s 46433 2181 46531 2279 4 gnd
port 3 nsew
rlabel metal3 s 42579 2950 42677 3048 4 gnd
port 3 nsew
rlabel metal3 s 43822 1979 43920 2077 4 gnd
port 3 nsew
rlabel metal3 s 49176 7426 49274 7524 4 gnd
port 3 nsew
rlabel metal3 s 45064 2513 45162 2611 4 vdd
port 2 nsew
rlabel metal3 s 43836 1563 43934 1661 4 vdd
port 2 nsew
rlabel metal3 s 42693 3743 42791 3841 4 gnd
port 3 nsew
rlabel metal3 s 42568 2513 42666 2611 4 vdd
port 2 nsew
rlabel metal3 s 46437 4065 46535 4163 4 vdd
port 2 nsew
rlabel metal3 s 42763 5677 42861 5775 4 gnd
port 3 nsew
rlabel metal3 s 46437 3743 46535 3841 4 gnd
port 3 nsew
rlabel metal3 s 42689 2181 42787 2279 4 gnd
port 3 nsew
rlabel metal3 s 46312 2513 46410 2611 4 vdd
port 2 nsew
rlabel metal3 s 46332 1563 46430 1661 4 vdd
port 2 nsew
rlabel metal3 s 45432 7426 45530 7524 4 gnd
port 3 nsew
rlabel metal3 s 47560 2513 47658 2611 4 vdd
port 2 nsew
rlabel metal3 s 43941 4065 44039 4163 4 vdd
port 2 nsew
rlabel metal3 s 46323 2950 46421 3048 4 gnd
port 3 nsew
rlabel metal3 s 42574 1979 42672 2077 4 gnd
port 3 nsew
rlabel metal3 s 48933 4065 49031 4163 4 vdd
port 2 nsew
rlabel metal3 s 46425 4903 46523 5001 4 vdd
port 2 nsew
rlabel metal3 s 48921 4903 49019 5001 4 vdd
port 2 nsew
rlabel metal3 s 47755 5677 47853 5775 4 gnd
port 3 nsew
rlabel metal3 s 45070 1979 45168 2077 4 gnd
port 3 nsew
rlabel metal3 s 49003 5677 49101 5775 4 gnd
port 3 nsew
rlabel metal3 s 43941 3743 44039 3841 4 gnd
port 3 nsew
rlabel metal3 s 45084 1563 45182 1661 4 vdd
port 2 nsew
rlabel metal3 s 47681 2181 47779 2279 4 gnd
port 3 nsew
rlabel metal3 s 47571 2950 47669 3048 4 gnd
port 3 nsew
rlabel metal3 s 44184 7426 44282 7524 4 gnd
port 3 nsew
rlabel metal3 s 43929 4903 44027 5001 4 vdd
port 2 nsew
rlabel metal3 s 42588 1563 42686 1661 4 vdd
port 2 nsew
rlabel metal3 s 46680 7426 46778 7524 4 gnd
port 3 nsew
rlabel metal3 s 48933 3743 49031 3841 4 gnd
port 3 nsew
rlabel metal3 s 41688 7426 41786 7524 4 gnd
port 3 nsew
rlabel metal3 s 42936 7426 43034 7524 4 gnd
port 3 nsew
rlabel metal3 s 64541 15285 64639 15383 4 gnd
port 3 nsew
rlabel metal3 s 65600 15262 65698 15360 4 vdd
port 2 nsew
rlabel metal3 s 63684 16075 63782 16173 4 vdd
port 2 nsew
rlabel metal3 s 63302 12892 63400 12990 4 gnd
port 3 nsew
rlabel metal3 s 63681 13689 63779 13787 4 vdd
port 2 nsew
rlabel metal3 s 64106 12899 64204 12997 4 gnd
port 3 nsew
rlabel metal3 s 62906 12892 63004 12990 4 vdd
port 2 nsew
rlabel metal3 s 65996 15262 66094 15360 4 gnd
port 3 nsew
rlabel metal3 s 63302 15262 63400 15360 4 gnd
port 3 nsew
rlabel metal3 s 65004 12892 65102 12990 4 vdd
port 2 nsew
rlabel metal3 s 64116 16075 64214 16173 4 vdd
port 2 nsew
rlabel metal3 s 64541 16075 64639 16173 4 gnd
port 3 nsew
rlabel metal3 s 63684 15285 63782 15383 4 vdd
port 2 nsew
rlabel metal3 s 63302 16052 63400 16150 4 gnd
port 3 nsew
rlabel metal3 s 62906 15262 63004 15360 4 vdd
port 2 nsew
rlabel metal3 s 64106 13689 64204 13787 4 gnd
port 3 nsew
rlabel metal3 s 64116 15285 64214 15383 4 vdd
port 2 nsew
rlabel metal3 s 62906 13682 63004 13780 4 vdd
port 2 nsew
rlabel metal3 s 65400 12892 65498 12990 4 gnd
port 3 nsew
rlabel metal3 s 62906 16052 63004 16150 4 vdd
port 2 nsew
rlabel metal3 s 63681 12899 63779 12997 4 vdd
port 2 nsew
rlabel metal3 s 63302 13682 63400 13780 4 gnd
port 3 nsew
rlabel metal3 s 60702 13705 60800 13803 4 vdd
port 2 nsew
rlabel metal3 s 59888 16052 59986 16150 4 gnd
port 3 nsew
rlabel metal3 s 61127 13331 61225 13429 4 gnd
port 3 nsew
rlabel metal3 s 61127 15701 61225 15799 4 gnd
port 3 nsew
rlabel metal3 s 60702 14853 60800 14951 4 vdd
port 2 nsew
rlabel metal3 s 61127 16075 61225 16173 4 gnd
port 3 nsew
rlabel metal3 s 60270 16075 60368 16173 4 vdd
port 2 nsew
rlabel metal3 s 61127 14121 61225 14219 4 gnd
port 3 nsew
rlabel metal3 s 59492 14472 59590 14570 4 vdd
port 2 nsew
rlabel metal3 s 61127 14911 61225 15009 4 gnd
port 3 nsew
rlabel metal3 s 60702 13273 60800 13371 4 vdd
port 2 nsew
rlabel metal3 s 60270 14495 60368 14593 4 vdd
port 2 nsew
rlabel metal3 s 60702 15643 60800 15741 4 vdd
port 2 nsew
rlabel metal3 s 60270 12915 60368 13013 4 vdd
port 2 nsew
rlabel metal3 s 59492 16052 59590 16150 4 vdd
port 2 nsew
rlabel metal3 s 60270 13273 60368 13371 4 vdd
port 2 nsew
rlabel metal3 s 59888 12892 59986 12990 4 gnd
port 3 nsew
rlabel metal3 s 59888 13682 59986 13780 4 gnd
port 3 nsew
rlabel metal3 s 60270 15285 60368 15383 4 vdd
port 2 nsew
rlabel metal3 s 59888 14472 59986 14570 4 gnd
port 3 nsew
rlabel metal3 s 59888 13287 59986 13385 4 gnd
port 3 nsew
rlabel metal3 s 61127 12915 61225 13013 4 gnd
port 3 nsew
rlabel metal3 s 61127 16491 61225 16589 4 gnd
port 3 nsew
rlabel metal3 s 60270 14063 60368 14161 4 vdd
port 2 nsew
rlabel metal3 s 59492 14077 59590 14175 4 vdd
port 2 nsew
rlabel metal3 s 60702 15285 60800 15383 4 vdd
port 2 nsew
rlabel metal3 s 60270 13705 60368 13803 4 vdd
port 2 nsew
rlabel metal3 s 59492 15657 59590 15755 4 vdd
port 2 nsew
rlabel metal3 s 59492 14867 59590 14965 4 vdd
port 2 nsew
rlabel metal3 s 61127 15285 61225 15383 4 gnd
port 3 nsew
rlabel metal3 s 60270 14853 60368 14951 4 vdd
port 2 nsew
rlabel metal3 s 59888 16447 59986 16545 4 gnd
port 3 nsew
rlabel metal3 s 59888 15262 59986 15360 4 gnd
port 3 nsew
rlabel metal3 s 60702 14063 60800 14161 4 vdd
port 2 nsew
rlabel metal3 s 60702 12915 60800 13013 4 vdd
port 2 nsew
rlabel metal3 s 59492 16447 59590 16545 4 vdd
port 2 nsew
rlabel metal3 s 61127 14495 61225 14593 4 gnd
port 3 nsew
rlabel metal3 s 60702 14495 60800 14593 4 vdd
port 2 nsew
rlabel metal3 s 59492 13682 59590 13780 4 vdd
port 2 nsew
rlabel metal3 s 61127 13705 61225 13803 4 gnd
port 3 nsew
rlabel metal3 s 59888 15657 59986 15755 4 gnd
port 3 nsew
rlabel metal3 s 60702 16075 60800 16173 4 vdd
port 2 nsew
rlabel metal3 s 59492 13287 59590 13385 4 vdd
port 2 nsew
rlabel metal3 s 59492 15262 59590 15360 4 vdd
port 2 nsew
rlabel metal3 s 59492 12892 59590 12990 4 vdd
port 2 nsew
rlabel metal3 s 60270 16433 60368 16531 4 vdd
port 2 nsew
rlabel metal3 s 59888 14077 59986 14175 4 gnd
port 3 nsew
rlabel metal3 s 60270 15643 60368 15741 4 vdd
port 2 nsew
rlabel metal3 s 59888 14867 59986 14965 4 gnd
port 3 nsew
rlabel metal3 s 60702 16433 60800 16531 4 vdd
port 2 nsew
rlabel metal3 s 60270 10903 60368 11001 4 vdd
port 2 nsew
rlabel metal3 s 61127 12541 61225 12639 4 gnd
port 3 nsew
rlabel metal3 s 61127 10545 61225 10643 4 gnd
port 3 nsew
rlabel metal3 s 60270 11693 60368 11791 4 vdd
port 2 nsew
rlabel metal3 s 60702 12125 60800 12223 4 vdd
port 2 nsew
rlabel metal3 s 59492 10917 59590 11015 4 vdd
port 2 nsew
rlabel metal3 s 60702 11693 60800 11791 4 vdd
port 2 nsew
rlabel metal3 s 61127 11335 61225 11433 4 gnd
port 3 nsew
rlabel metal3 s 60270 11335 60368 11433 4 vdd
port 2 nsew
rlabel metal3 s 60702 11335 60800 11433 4 vdd
port 2 nsew
rlabel metal3 s 59888 10522 59986 10620 4 gnd
port 3 nsew
rlabel metal3 s 60270 12483 60368 12581 4 vdd
port 2 nsew
rlabel metal3 s 60270 12125 60368 12223 4 vdd
port 2 nsew
rlabel metal3 s 61127 10961 61225 11059 4 gnd
port 3 nsew
rlabel metal3 s 59888 12102 59986 12200 4 gnd
port 3 nsew
rlabel metal3 s 59492 12497 59590 12595 4 vdd
port 2 nsew
rlabel metal3 s 61127 12125 61225 12223 4 gnd
port 3 nsew
rlabel metal3 s 60702 12483 60800 12581 4 vdd
port 2 nsew
rlabel metal3 s 60702 10903 60800 11001 4 vdd
port 2 nsew
rlabel metal3 s 59888 10917 59986 11015 4 gnd
port 3 nsew
rlabel metal3 s 59888 12497 59986 12595 4 gnd
port 3 nsew
rlabel metal3 s 59888 11312 59986 11410 4 gnd
port 3 nsew
rlabel metal3 s 59492 11312 59590 11410 4 vdd
port 2 nsew
rlabel metal3 s 59492 10522 59590 10620 4 vdd
port 2 nsew
rlabel metal3 s 61127 11751 61225 11849 4 gnd
port 3 nsew
rlabel metal3 s 60702 10545 60800 10643 4 vdd
port 2 nsew
rlabel metal3 s 60270 10545 60368 10643 4 vdd
port 2 nsew
rlabel metal3 s 59492 11707 59590 11805 4 vdd
port 2 nsew
rlabel metal3 s 59888 11707 59986 11805 4 gnd
port 3 nsew
rlabel metal3 s 59492 12102 59590 12200 4 vdd
port 2 nsew
rlabel metal3 s 64106 10529 64204 10627 4 gnd
port 3 nsew
rlabel metal3 s 63302 11312 63400 11410 4 gnd
port 3 nsew
rlabel metal3 s 62906 10522 63004 10620 4 vdd
port 2 nsew
rlabel metal3 s 62906 11312 63004 11410 4 vdd
port 2 nsew
rlabel metal3 s 64106 11319 64204 11417 4 gnd
port 3 nsew
rlabel metal3 s 63302 10522 63400 10620 4 gnd
port 3 nsew
rlabel metal3 s 63681 10529 63779 10627 4 vdd
port 2 nsew
rlabel metal3 s 63681 11319 63779 11417 4 vdd
port 2 nsew
rlabel metal3 s 65400 10522 65498 10620 4 gnd
port 3 nsew
rlabel metal3 s 65004 10522 65102 10620 4 vdd
port 2 nsew
rlabel metal3 s 54552 11154 54650 11252 4 gnd
port 3 nsew
rlabel metal3 s 54552 10917 54650 11015 4 gnd
port 3 nsew
rlabel metal3 s 51241 8975 51339 9073 4 vdd
port 2 nsew
rlabel metal3 s 54552 15104 54650 15202 4 gnd
port 3 nsew
rlabel metal3 s 54552 13287 54650 13385 4 gnd
port 3 nsew
rlabel metal3 s 54552 12260 54650 12358 4 gnd
port 3 nsew
rlabel metal3 s 54552 10127 54650 10225 4 gnd
port 3 nsew
rlabel metal3 s 54552 14867 54650 14965 4 gnd
port 3 nsew
rlabel metal3 s 50112 9566 50210 9664 4 vdd
port 2 nsew
rlabel metal3 s 52103 8975 52201 9073 4 vdd
port 2 nsew
rlabel metal3 s 54552 12497 54650 12595 4 gnd
port 3 nsew
rlabel metal3 s 54552 13524 54650 13622 4 gnd
port 3 nsew
rlabel metal3 s 54552 16447 54650 16545 4 gnd
port 3 nsew
rlabel metal3 s 50736 9566 50834 9664 4 vdd
port 2 nsew
rlabel metal3 s 54918 10000 55016 10098 4 gnd
port 3 nsew
rlabel metal3 s 53351 8975 53449 9073 4 vdd
port 2 nsew
rlabel metal3 s 54552 10364 54650 10462 4 gnd
port 3 nsew
rlabel metal3 s 52608 9566 52706 9664 4 vdd
port 2 nsew
rlabel metal3 s 53232 9566 53330 9664 4 vdd
port 2 nsew
rlabel metal3 s 53856 9566 53954 9664 4 vdd
port 2 nsew
rlabel metal3 s 54552 11470 54650 11568 4 gnd
port 3 nsew
rlabel metal3 s 54552 15657 54650 15755 4 gnd
port 3 nsew
rlabel metal3 s 54552 14077 54650 14175 4 gnd
port 3 nsew
rlabel metal3 s 50855 8975 50953 9073 4 vdd
port 2 nsew
rlabel metal3 s 51360 9566 51458 9664 4 vdd
port 2 nsew
rlabel metal3 s 54552 11707 54650 11805 4 gnd
port 3 nsew
rlabel metal3 s 54552 13840 54650 13938 4 gnd
port 3 nsew
rlabel metal3 s 54552 13050 54650 13148 4 gnd
port 3 nsew
rlabel metal3 s 51984 9566 52082 9664 4 vdd
port 2 nsew
rlabel metal3 s 54552 11944 54650 12042 4 gnd
port 3 nsew
rlabel metal3 s 54552 14314 54650 14412 4 gnd
port 3 nsew
rlabel metal3 s 54552 10680 54650 10778 4 gnd
port 3 nsew
rlabel metal3 s 52489 8975 52587 9073 4 vdd
port 2 nsew
rlabel metal3 s 49993 8975 50091 9073 4 vdd
port 2 nsew
rlabel metal3 s 54552 16210 54650 16308 4 gnd
port 3 nsew
rlabel metal3 s 54552 15420 54650 15518 4 gnd
port 3 nsew
rlabel metal3 s 54552 12734 54650 12832 4 gnd
port 3 nsew
rlabel metal3 s 54552 14630 54650 14728 4 gnd
port 3 nsew
rlabel metal3 s 54552 16684 54650 16782 4 gnd
port 3 nsew
rlabel metal3 s 54552 15894 54650 15992 4 gnd
port 3 nsew
rlabel metal3 s 50076 1563 50174 1661 4 vdd
port 2 nsew
rlabel metal3 s 51672 7426 51770 7524 4 gnd
port 3 nsew
rlabel metal3 s 50169 4903 50267 5001 4 vdd
port 2 nsew
rlabel metal3 s 51304 2513 51402 2611 4 vdd
port 2 nsew
rlabel metal3 s 52677 3743 52775 3841 4 gnd
port 3 nsew
rlabel metal3 s 50062 1979 50160 2077 4 gnd
port 3 nsew
rlabel metal3 s 51324 1563 51422 1661 4 vdd
port 2 nsew
rlabel metal3 s 50251 5677 50349 5775 4 gnd
port 3 nsew
rlabel metal3 s 52920 7426 53018 7524 4 gnd
port 3 nsew
rlabel metal3 s 51417 4903 51515 5001 4 vdd
port 2 nsew
rlabel metal3 s 51499 5677 51597 5775 4 gnd
port 3 nsew
rlabel metal3 s 52673 2181 52771 2279 4 gnd
port 3 nsew
rlabel metal3 s 50181 4065 50279 4163 4 vdd
port 2 nsew
rlabel metal3 s 52747 5677 52845 5775 4 gnd
port 3 nsew
rlabel metal3 s 53544 1120 53642 1218 4 vdd
port 2 nsew
rlabel metal3 s 50177 2181 50275 2279 4 gnd
port 3 nsew
rlabel metal3 s 51425 2181 51523 2279 4 gnd
port 3 nsew
rlabel metal3 s 52552 2513 52650 2611 4 vdd
port 2 nsew
rlabel metal3 s 51429 4065 51527 4163 4 vdd
port 2 nsew
rlabel metal3 s 50056 2513 50154 2611 4 vdd
port 2 nsew
rlabel metal3 s 52677 4065 52775 4163 4 vdd
port 2 nsew
rlabel metal3 s 51429 3743 51527 3841 4 gnd
port 3 nsew
rlabel metal3 s 52563 2950 52661 3048 4 gnd
port 3 nsew
rlabel metal3 s 51310 1979 51408 2077 4 gnd
port 3 nsew
rlabel metal3 s 50424 7426 50522 7524 4 gnd
port 3 nsew
rlabel metal3 s 51315 2950 51413 3048 4 gnd
port 3 nsew
rlabel metal3 s 50067 2950 50165 3048 4 gnd
port 3 nsew
rlabel metal3 s 52572 1563 52670 1661 4 vdd
port 2 nsew
rlabel metal3 s 50181 3743 50279 3841 4 gnd
port 3 nsew
rlabel metal3 s 52558 1979 52656 2077 4 gnd
port 3 nsew
rlabel metal3 s 53544 0 53642 98 4 gnd
port 3 nsew
rlabel metal3 s 52665 4903 52763 5001 4 vdd
port 2 nsew
rlabel metal2 s 11663 49 11691 9386 4 p_en_bar0
port 5 nsew
rlabel metal2 s 11787 49 11815 9386 4 s_en0
port 6 nsew
rlabel metal2 s 11911 49 11939 9386 4 w_en0
port 7 nsew
rlabel metal2 s 7960 9863 7988 9891 4 wl_en0
port 8 nsew
rlabel metal2 s 55277 61526 55305 67312 4 s_en1
port 9 nsew
rlabel metal2 s 55401 61526 55429 67312 4 p_en_bar1
port 10 nsew
rlabel metal2 s 59262 61021 59290 61049 4 wl_en1
port 11 nsew
rlabel metal2 s 13643 305 13671 333 4 bank_wmask0_0
port 12 nsew
rlabel metal2 s 23627 305 23655 333 4 bank_wmask0_1
port 13 nsew
rlabel metal2 s 33611 305 33639 333 4 bank_wmask0_2
port 14 nsew
rlabel metal2 s 43595 305 43623 333 4 bank_wmask0_3
port 15 nsew
rlabel metal1 s 33729 66974 33775 67228 4 dout1_16
port 16 nsew
rlabel metal1 s 34977 66974 35023 67228 4 dout1_17
port 17 nsew
rlabel metal1 s 36225 66974 36271 67228 4 dout1_18
port 18 nsew
rlabel metal1 s 37473 66974 37519 67228 4 dout1_19
port 19 nsew
rlabel metal1 s 38721 66974 38767 67228 4 dout1_20
port 20 nsew
rlabel metal1 s 39969 66974 40015 67228 4 dout1_21
port 21 nsew
rlabel metal1 s 41217 66974 41263 67228 4 dout1_22
port 22 nsew
rlabel metal1 s 42465 66974 42511 67228 4 dout1_23
port 23 nsew
rlabel metal1 s 43713 66974 43759 67228 4 dout1_24
port 24 nsew
rlabel metal1 s 44961 66974 45007 67228 4 dout1_25
port 25 nsew
rlabel metal1 s 46209 66974 46255 67228 4 dout1_26
port 26 nsew
rlabel metal1 s 47457 66974 47503 67228 4 dout1_27
port 27 nsew
rlabel metal1 s 48705 66974 48751 67228 4 dout1_28
port 28 nsew
rlabel metal1 s 49953 66974 49999 67228 4 dout1_29
port 29 nsew
rlabel metal1 s 51201 66974 51247 67228 4 dout1_30
port 30 nsew
rlabel metal1 s 52449 66974 52495 67228 4 dout1_31
port 31 nsew
rlabel metal1 s 13761 66974 13807 67228 4 dout1_0
port 32 nsew
rlabel metal1 s 15009 66974 15055 67228 4 dout1_1
port 33 nsew
rlabel metal1 s 16257 66974 16303 67228 4 dout1_2
port 34 nsew
rlabel metal1 s 17505 66974 17551 67228 4 dout1_3
port 35 nsew
rlabel metal1 s 18753 66974 18799 67228 4 dout1_4
port 36 nsew
rlabel metal1 s 20001 66974 20047 67228 4 dout1_5
port 37 nsew
rlabel metal1 s 21249 66974 21295 67228 4 dout1_6
port 38 nsew
rlabel metal1 s 22497 66974 22543 67228 4 dout1_7
port 39 nsew
rlabel metal1 s 23745 66974 23791 67228 4 dout1_8
port 40 nsew
rlabel metal1 s 24993 66974 25039 67228 4 dout1_9
port 41 nsew
rlabel metal1 s 26241 66974 26287 67228 4 dout1_10
port 42 nsew
rlabel metal1 s 27489 66974 27535 67228 4 dout1_11
port 43 nsew
rlabel metal1 s 28737 66974 28783 67228 4 dout1_12
port 44 nsew
rlabel metal1 s 29985 66974 30031 67228 4 dout1_13
port 45 nsew
rlabel metal1 s 31233 66974 31279 67228 4 dout1_14
port 46 nsew
rlabel metal1 s 32481 66974 32527 67228 4 dout1_15
port 47 nsew
rlabel metal1 s 19 10176 47 18076 4 addr0_1
port 48 nsew
rlabel metal1 s 99 10176 127 18076 4 addr0_2
port 49 nsew
rlabel metal1 s 179 10176 207 18076 4 addr0_3
port 50 nsew
rlabel metal1 s 259 10176 287 18076 4 addr0_4
port 51 nsew
rlabel metal1 s 339 10176 367 18076 4 addr0_5
port 52 nsew
rlabel metal1 s 419 10176 447 18076 4 addr0_6
port 53 nsew
rlabel metal1 s 499 10176 527 18076 4 addr0_7
port 54 nsew
rlabel metal1 s 13912 1425 13972 1481 4 din0_0
port 55 nsew
rlabel metal1 s 15160 1425 15220 1481 4 din0_1
port 56 nsew
rlabel metal1 s 16408 1425 16468 1481 4 din0_2
port 57 nsew
rlabel metal1 s 17656 1425 17716 1481 4 din0_3
port 58 nsew
rlabel metal1 s 18904 1425 18964 1481 4 din0_4
port 59 nsew
rlabel metal1 s 20152 1425 20212 1481 4 din0_5
port 60 nsew
rlabel metal1 s 21400 1425 21460 1481 4 din0_6
port 61 nsew
rlabel metal1 s 22648 1425 22708 1481 4 din0_7
port 62 nsew
rlabel metal1 s 23896 1425 23956 1481 4 din0_8
port 63 nsew
rlabel metal1 s 25144 1425 25204 1481 4 din0_9
port 64 nsew
rlabel metal1 s 26392 1425 26452 1481 4 din0_10
port 65 nsew
rlabel metal1 s 27640 1425 27700 1481 4 din0_11
port 66 nsew
rlabel metal1 s 28888 1425 28948 1481 4 din0_12
port 67 nsew
rlabel metal1 s 30136 1425 30196 1481 4 din0_13
port 68 nsew
rlabel metal1 s 31384 1425 31444 1481 4 din0_14
port 69 nsew
rlabel metal1 s 32632 1425 32692 1481 4 din0_15
port 70 nsew
rlabel metal1 s 13761 3684 13807 3938 4 dout0_0
port 71 nsew
rlabel metal1 s 15009 3684 15055 3938 4 dout0_1
port 72 nsew
rlabel metal1 s 16257 3684 16303 3938 4 dout0_2
port 73 nsew
rlabel metal1 s 17505 3684 17551 3938 4 dout0_3
port 74 nsew
rlabel metal1 s 18753 3684 18799 3938 4 dout0_4
port 75 nsew
rlabel metal1 s 20001 3684 20047 3938 4 dout0_5
port 76 nsew
rlabel metal1 s 21249 3684 21295 3938 4 dout0_6
port 77 nsew
rlabel metal1 s 22497 3684 22543 3938 4 dout0_7
port 78 nsew
rlabel metal1 s 23745 3684 23791 3938 4 dout0_8
port 79 nsew
rlabel metal1 s 24993 3684 25039 3938 4 dout0_9
port 80 nsew
rlabel metal1 s 26241 3684 26287 3938 4 dout0_10
port 81 nsew
rlabel metal1 s 27489 3684 27535 3938 4 dout0_11
port 82 nsew
rlabel metal1 s 28737 3684 28783 3938 4 dout0_12
port 83 nsew
rlabel metal1 s 29985 3684 30031 3938 4 dout0_13
port 84 nsew
rlabel metal1 s 31233 3684 31279 3938 4 dout0_14
port 85 nsew
rlabel metal1 s 32481 3684 32527 3938 4 dout0_15
port 86 nsew
rlabel metal1 s 42616 1425 42676 1481 4 din0_23
port 87 nsew
rlabel metal1 s 43864 1425 43924 1481 4 din0_24
port 88 nsew
rlabel metal1 s 45112 1425 45172 1481 4 din0_25
port 89 nsew
rlabel metal1 s 46360 1425 46420 1481 4 din0_26
port 90 nsew
rlabel metal1 s 47608 1425 47668 1481 4 din0_27
port 91 nsew
rlabel metal1 s 48856 1425 48916 1481 4 din0_28
port 92 nsew
rlabel metal1 s 50104 1425 50164 1481 4 din0_29
port 93 nsew
rlabel metal1 s 51352 1425 51412 1481 4 din0_30
port 94 nsew
rlabel metal1 s 52600 1425 52660 1481 4 din0_31
port 95 nsew
rlabel metal1 s 33729 3684 33775 3938 4 dout0_16
port 96 nsew
rlabel metal1 s 34977 3684 35023 3938 4 dout0_17
port 97 nsew
rlabel metal1 s 36225 3684 36271 3938 4 dout0_18
port 98 nsew
rlabel metal1 s 37473 3684 37519 3938 4 dout0_19
port 99 nsew
rlabel metal1 s 38721 3684 38767 3938 4 dout0_20
port 100 nsew
rlabel metal1 s 39969 3684 40015 3938 4 dout0_21
port 101 nsew
rlabel metal1 s 41217 3684 41263 3938 4 dout0_22
port 102 nsew
rlabel metal1 s 42465 3684 42511 3938 4 dout0_23
port 103 nsew
rlabel metal1 s 43713 3684 43759 3938 4 dout0_24
port 104 nsew
rlabel metal1 s 44961 3684 45007 3938 4 dout0_25
port 105 nsew
rlabel metal1 s 46209 3684 46255 3938 4 dout0_26
port 106 nsew
rlabel metal1 s 47457 3684 47503 3938 4 dout0_27
port 107 nsew
rlabel metal1 s 48705 3684 48751 3938 4 dout0_28
port 108 nsew
rlabel metal1 s 49953 3684 49999 3938 4 dout0_29
port 109 nsew
rlabel metal1 s 51201 3684 51247 3938 4 dout0_30
port 110 nsew
rlabel metal1 s 52449 3684 52495 3938 4 dout0_31
port 111 nsew
rlabel metal1 s 33880 1425 33940 1481 4 din0_16
port 112 nsew
rlabel metal1 s 35128 1425 35188 1481 4 din0_17
port 113 nsew
rlabel metal1 s 36376 1425 36436 1481 4 din0_18
port 114 nsew
rlabel metal1 s 37624 1425 37684 1481 4 din0_19
port 115 nsew
rlabel metal1 s 38872 1425 38932 1481 4 din0_20
port 116 nsew
rlabel metal1 s 40120 1425 40180 1481 4 din0_21
port 117 nsew
rlabel metal1 s 41368 1425 41428 1481 4 din0_22
port 118 nsew
rlabel metal1 s 67203 10176 67231 18076 4 addr1_1
port 119 nsew
rlabel metal1 s 67123 10176 67151 18076 4 addr1_2
port 120 nsew
rlabel metal1 s 67043 10176 67071 18076 4 addr1_3
port 121 nsew
rlabel metal1 s 66963 10176 66991 18076 4 addr1_4
port 122 nsew
rlabel metal1 s 66883 10176 66911 18076 4 addr1_5
port 123 nsew
rlabel metal1 s 66803 10176 66831 18076 4 addr1_6
port 124 nsew
rlabel metal1 s 66723 10176 66751 18076 4 addr1_7
port 125 nsew
rlabel locali s 6070 5476 6070 5476 4 addr0_0
port 126 nsew
rlabel locali s 61056 65436 61056 65436 4 addr1_0
port 127 nsew
<< properties >>
string FIXED_BBOX 0 0 67334 67263
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_END 8110094
string GDS_START 7440238
<< end >>
