(* blackbox *)
module scs8hvl_lsbufhv2lv_1(input A, output X); endmodule   
(* blackbox *)
module scs8hvl_lsbuflv2hv_1(input A, output X); endmodule   
