magic
tech sky130A
magscale 1 2
timestamp 1636140361
<< checkpaint >>
rect -1319 -1316 2873 1714
<< nwell >>
rect -54 284 1608 454
rect -59 116 1613 284
rect -54 -54 1608 116
<< scpmos >>
rect 60 0 90 400
rect 168 0 198 400
rect 276 0 306 400
rect 384 0 414 400
rect 492 0 522 400
rect 600 0 630 400
rect 708 0 738 400
rect 816 0 846 400
rect 924 0 954 400
rect 1032 0 1062 400
rect 1140 0 1170 400
rect 1248 0 1278 400
rect 1356 0 1386 400
rect 1464 0 1494 400
<< pdiff >>
rect 0 217 60 400
rect 0 183 8 217
rect 42 183 60 217
rect 0 0 60 183
rect 90 217 168 400
rect 90 183 112 217
rect 146 183 168 217
rect 90 0 168 183
rect 198 217 276 400
rect 198 183 220 217
rect 254 183 276 217
rect 198 0 276 183
rect 306 217 384 400
rect 306 183 328 217
rect 362 183 384 217
rect 306 0 384 183
rect 414 217 492 400
rect 414 183 436 217
rect 470 183 492 217
rect 414 0 492 183
rect 522 217 600 400
rect 522 183 544 217
rect 578 183 600 217
rect 522 0 600 183
rect 630 217 708 400
rect 630 183 652 217
rect 686 183 708 217
rect 630 0 708 183
rect 738 217 816 400
rect 738 183 760 217
rect 794 183 816 217
rect 738 0 816 183
rect 846 217 924 400
rect 846 183 868 217
rect 902 183 924 217
rect 846 0 924 183
rect 954 217 1032 400
rect 954 183 976 217
rect 1010 183 1032 217
rect 954 0 1032 183
rect 1062 217 1140 400
rect 1062 183 1084 217
rect 1118 183 1140 217
rect 1062 0 1140 183
rect 1170 217 1248 400
rect 1170 183 1192 217
rect 1226 183 1248 217
rect 1170 0 1248 183
rect 1278 217 1356 400
rect 1278 183 1300 217
rect 1334 183 1356 217
rect 1278 0 1356 183
rect 1386 217 1464 400
rect 1386 183 1408 217
rect 1442 183 1464 217
rect 1386 0 1464 183
rect 1494 217 1554 400
rect 1494 183 1512 217
rect 1546 183 1554 217
rect 1494 0 1554 183
<< pdiffc >>
rect 8 183 42 217
rect 112 183 146 217
rect 220 183 254 217
rect 328 183 362 217
rect 436 183 470 217
rect 544 183 578 217
rect 652 183 686 217
rect 760 183 794 217
rect 868 183 902 217
rect 976 183 1010 217
rect 1084 183 1118 217
rect 1192 183 1226 217
rect 1300 183 1334 217
rect 1408 183 1442 217
rect 1512 183 1546 217
<< poly >>
rect 60 400 90 426
rect 168 400 198 426
rect 276 400 306 426
rect 384 400 414 426
rect 492 400 522 426
rect 600 400 630 426
rect 708 400 738 426
rect 816 400 846 426
rect 924 400 954 426
rect 1032 400 1062 426
rect 1140 400 1170 426
rect 1248 400 1278 426
rect 1356 400 1386 426
rect 1464 400 1494 426
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 1356 -26 1386 0
rect 1464 -26 1494 0
rect 60 -56 1494 -26
<< locali >>
rect 8 217 42 233
rect 8 167 42 183
rect 112 217 146 233
rect 112 133 146 183
rect 220 217 254 233
rect 220 167 254 183
rect 328 217 362 233
rect 328 133 362 183
rect 436 217 470 233
rect 436 167 470 183
rect 544 217 578 233
rect 544 133 578 183
rect 652 217 686 233
rect 652 167 686 183
rect 760 217 794 233
rect 760 133 794 183
rect 868 217 902 233
rect 868 167 902 183
rect 976 217 1010 233
rect 976 133 1010 183
rect 1084 217 1118 233
rect 1084 167 1118 183
rect 1192 217 1226 233
rect 1192 133 1226 183
rect 1300 217 1334 233
rect 1300 167 1334 183
rect 1408 217 1442 233
rect 1408 133 1442 183
rect 1512 217 1546 233
rect 1512 167 1546 183
rect 112 99 1442 133
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_0
timestamp 1636140361
transform 1 0 1504 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_1
timestamp 1636140361
transform 1 0 1400 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_2
timestamp 1636140361
transform 1 0 1292 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_3
timestamp 1636140361
transform 1 0 1184 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_4
timestamp 1636140361
transform 1 0 1076 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_5
timestamp 1636140361
transform 1 0 968 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_6
timestamp 1636140361
transform 1 0 860 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_7
timestamp 1636140361
transform 1 0 752 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_8
timestamp 1636140361
transform 1 0 644 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_9
timestamp 1636140361
transform 1 0 536 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_10
timestamp 1636140361
transform 1 0 428 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_11
timestamp 1636140361
transform 1 0 320 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_12
timestamp 1636140361
transform 1 0 212 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_13
timestamp 1636140361
transform 1 0 104 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_14
timestamp 1636140361
transform 1 0 0 0 1 167
box 0 0 1 1
<< labels >>
rlabel locali s 453 200 453 200 4 S
port 1 nsew
rlabel locali s 1529 200 1529 200 4 S
port 1 nsew
rlabel locali s 25 200 25 200 4 S
port 1 nsew
rlabel locali s 885 200 885 200 4 S
port 1 nsew
rlabel locali s 1317 200 1317 200 4 S
port 1 nsew
rlabel locali s 1101 200 1101 200 4 S
port 1 nsew
rlabel locali s 237 200 237 200 4 S
port 1 nsew
rlabel locali s 669 200 669 200 4 S
port 1 nsew
rlabel locali s 777 116 777 116 4 D
port 2 nsew
rlabel poly s 777 -41 777 -41 4 G
port 3 nsew
<< properties >>
string FIXED_BBOX -54 -56 1608 116
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_END 97864
string GDS_START 94006
<< end >>
