magic
tech sky130A
magscale 1 2
timestamp 1636140361
<< checkpaint >>
rect -1296 -1309 3136 11397
<< locali >>
rect 639 10097 673 10113
rect 639 10047 673 10063
rect 1375 10097 1409 10113
rect 1375 10047 1409 10063
rect 64 9499 98 9515
rect 64 9449 98 9465
rect 179 9499 213 9515
rect 179 9449 213 9465
rect 432 9499 466 9515
rect 432 9449 466 9465
rect 800 9499 834 9515
rect 800 9449 834 9465
rect 1168 9499 1202 9515
rect 1168 9449 1202 9465
rect 1536 9499 1570 9515
rect 1536 9449 1570 9465
rect 639 8977 673 8993
rect 639 8927 673 8943
rect 1375 8977 1409 8993
rect 1375 8927 1409 8943
rect 64 8455 98 8471
rect 64 8405 98 8421
rect 179 8455 213 8471
rect 179 8405 213 8421
rect 432 8455 466 8471
rect 432 8405 466 8421
rect 800 8455 834 8471
rect 800 8405 834 8421
rect 1168 8455 1202 8471
rect 1168 8405 1202 8421
rect 1536 8455 1570 8471
rect 1536 8405 1570 8421
rect 639 7857 673 7873
rect 639 7807 673 7823
rect 1375 7857 1409 7873
rect 1375 7807 1409 7823
rect 64 7259 98 7275
rect 64 7209 98 7225
rect 179 7259 213 7275
rect 179 7209 213 7225
rect 432 7259 466 7275
rect 432 7209 466 7225
rect 800 7259 834 7275
rect 800 7209 834 7225
rect 1168 7259 1202 7275
rect 1168 7209 1202 7225
rect 1536 7259 1570 7275
rect 1536 7209 1570 7225
rect 639 6737 673 6753
rect 639 6687 673 6703
rect 1375 6737 1409 6753
rect 1375 6687 1409 6703
rect 64 6215 98 6231
rect 64 6165 98 6181
rect 179 6215 213 6231
rect 179 6165 213 6181
rect 432 6215 466 6231
rect 432 6165 466 6181
rect 800 6215 834 6231
rect 800 6165 834 6181
rect 1168 6215 1202 6231
rect 1168 6165 1202 6181
rect 1536 6215 1570 6231
rect 1536 6165 1570 6181
rect 639 5617 673 5633
rect 639 5567 673 5583
rect 1375 5617 1409 5633
rect 1375 5567 1409 5583
rect 64 5019 98 5035
rect 64 4969 98 4985
rect 179 5019 213 5035
rect 179 4969 213 4985
rect 432 5019 466 5035
rect 432 4969 466 4985
rect 800 5019 834 5035
rect 800 4969 834 4985
rect 1168 5019 1202 5035
rect 1168 4969 1202 4985
rect 1536 5019 1570 5035
rect 1536 4969 1570 4985
rect 639 4497 673 4513
rect 639 4447 673 4463
rect 1375 4497 1409 4513
rect 1375 4447 1409 4463
rect 64 3975 98 3991
rect 64 3925 98 3941
rect 179 3975 213 3991
rect 179 3925 213 3941
rect 432 3975 466 3991
rect 432 3925 466 3941
rect 800 3975 834 3991
rect 800 3925 834 3941
rect 1168 3975 1202 3991
rect 1168 3925 1202 3941
rect 1536 3975 1570 3991
rect 1536 3925 1570 3941
rect 639 3377 673 3393
rect 639 3327 673 3343
rect 1375 3377 1409 3393
rect 1375 3327 1409 3343
rect 64 2779 98 2795
rect 64 2729 98 2745
rect 179 2779 213 2795
rect 179 2729 213 2745
rect 432 2779 466 2795
rect 432 2729 466 2745
rect 800 2779 834 2795
rect 800 2729 834 2745
rect 1168 2779 1202 2795
rect 1168 2729 1202 2745
rect 1536 2779 1570 2795
rect 1536 2729 1570 2745
rect 639 2257 673 2273
rect 639 2207 673 2223
rect 1375 2257 1409 2273
rect 1375 2207 1409 2223
rect 64 1735 98 1751
rect 64 1685 98 1701
rect 179 1735 213 1751
rect 179 1685 213 1701
rect 432 1735 466 1751
rect 432 1685 466 1701
rect 800 1735 834 1751
rect 800 1685 834 1701
rect 1168 1735 1202 1751
rect 1168 1685 1202 1701
rect 1536 1735 1570 1751
rect 1536 1685 1570 1701
rect 639 1137 673 1153
rect 639 1087 673 1103
rect 1375 1137 1409 1153
rect 1375 1087 1409 1103
rect 64 539 98 555
rect 64 489 98 505
rect 179 539 213 555
rect 179 489 213 505
rect 432 539 466 555
rect 432 489 466 505
rect 800 539 834 555
rect 800 489 834 505
rect 1168 539 1202 555
rect 1168 489 1202 505
rect 1536 539 1570 555
rect 1536 489 1570 505
rect 639 17 673 33
rect 639 -33 673 -17
rect 1375 17 1409 33
rect 1375 -33 1409 -17
<< viali >>
rect 639 10063 673 10097
rect 1375 10063 1409 10097
rect 64 9465 98 9499
rect 179 9465 213 9499
rect 432 9465 466 9499
rect 800 9465 834 9499
rect 1168 9465 1202 9499
rect 1536 9465 1570 9499
rect 639 8943 673 8977
rect 1375 8943 1409 8977
rect 64 8421 98 8455
rect 179 8421 213 8455
rect 432 8421 466 8455
rect 800 8421 834 8455
rect 1168 8421 1202 8455
rect 1536 8421 1570 8455
rect 639 7823 673 7857
rect 1375 7823 1409 7857
rect 64 7225 98 7259
rect 179 7225 213 7259
rect 432 7225 466 7259
rect 800 7225 834 7259
rect 1168 7225 1202 7259
rect 1536 7225 1570 7259
rect 639 6703 673 6737
rect 1375 6703 1409 6737
rect 64 6181 98 6215
rect 179 6181 213 6215
rect 432 6181 466 6215
rect 800 6181 834 6215
rect 1168 6181 1202 6215
rect 1536 6181 1570 6215
rect 639 5583 673 5617
rect 1375 5583 1409 5617
rect 64 4985 98 5019
rect 179 4985 213 5019
rect 432 4985 466 5019
rect 800 4985 834 5019
rect 1168 4985 1202 5019
rect 1536 4985 1570 5019
rect 639 4463 673 4497
rect 1375 4463 1409 4497
rect 64 3941 98 3975
rect 179 3941 213 3975
rect 432 3941 466 3975
rect 800 3941 834 3975
rect 1168 3941 1202 3975
rect 1536 3941 1570 3975
rect 639 3343 673 3377
rect 1375 3343 1409 3377
rect 64 2745 98 2779
rect 179 2745 213 2779
rect 432 2745 466 2779
rect 800 2745 834 2779
rect 1168 2745 1202 2779
rect 1536 2745 1570 2779
rect 639 2223 673 2257
rect 1375 2223 1409 2257
rect 64 1701 98 1735
rect 179 1701 213 1735
rect 432 1701 466 1735
rect 800 1701 834 1735
rect 1168 1701 1202 1735
rect 1536 1701 1570 1735
rect 639 1103 673 1137
rect 1375 1103 1409 1137
rect 64 505 98 539
rect 179 505 213 539
rect 432 505 466 539
rect 800 505 834 539
rect 1168 505 1202 539
rect 1536 505 1570 539
rect 639 -17 673 17
rect 1375 -17 1409 17
<< metal1 >>
rect 624 10054 630 10106
rect 682 10054 688 10106
rect 1360 10054 1366 10106
rect 1418 10054 1424 10106
rect 49 9456 55 9508
rect 107 9456 113 9508
rect 164 9456 170 9508
rect 222 9456 228 9508
rect 417 9456 423 9508
rect 475 9456 481 9508
rect 785 9456 791 9508
rect 843 9456 849 9508
rect 1153 9456 1159 9508
rect 1211 9456 1217 9508
rect 1521 9456 1527 9508
rect 1579 9456 1585 9508
rect 624 8934 630 8986
rect 682 8934 688 8986
rect 1360 8934 1366 8986
rect 1418 8934 1424 8986
rect 49 8412 55 8464
rect 107 8412 113 8464
rect 164 8412 170 8464
rect 222 8412 228 8464
rect 417 8412 423 8464
rect 475 8412 481 8464
rect 785 8412 791 8464
rect 843 8412 849 8464
rect 1153 8412 1159 8464
rect 1211 8412 1217 8464
rect 1521 8412 1527 8464
rect 1579 8412 1585 8464
rect 624 7814 630 7866
rect 682 7814 688 7866
rect 1360 7814 1366 7866
rect 1418 7814 1424 7866
rect 49 7216 55 7268
rect 107 7216 113 7268
rect 164 7216 170 7268
rect 222 7216 228 7268
rect 417 7216 423 7268
rect 475 7216 481 7268
rect 785 7216 791 7268
rect 843 7216 849 7268
rect 1153 7216 1159 7268
rect 1211 7216 1217 7268
rect 1521 7216 1527 7268
rect 1579 7216 1585 7268
rect 624 6694 630 6746
rect 682 6694 688 6746
rect 1360 6694 1366 6746
rect 1418 6694 1424 6746
rect 49 6172 55 6224
rect 107 6172 113 6224
rect 164 6172 170 6224
rect 222 6172 228 6224
rect 417 6172 423 6224
rect 475 6172 481 6224
rect 785 6172 791 6224
rect 843 6172 849 6224
rect 1153 6172 1159 6224
rect 1211 6172 1217 6224
rect 1521 6172 1527 6224
rect 1579 6172 1585 6224
rect 624 5574 630 5626
rect 682 5574 688 5626
rect 1360 5574 1366 5626
rect 1418 5574 1424 5626
rect 49 4976 55 5028
rect 107 4976 113 5028
rect 164 4976 170 5028
rect 222 4976 228 5028
rect 417 4976 423 5028
rect 475 4976 481 5028
rect 785 4976 791 5028
rect 843 4976 849 5028
rect 1153 4976 1159 5028
rect 1211 4976 1217 5028
rect 1521 4976 1527 5028
rect 1579 4976 1585 5028
rect 624 4454 630 4506
rect 682 4454 688 4506
rect 1360 4454 1366 4506
rect 1418 4454 1424 4506
rect 49 3932 55 3984
rect 107 3932 113 3984
rect 164 3932 170 3984
rect 222 3932 228 3984
rect 417 3932 423 3984
rect 475 3932 481 3984
rect 785 3932 791 3984
rect 843 3932 849 3984
rect 1153 3932 1159 3984
rect 1211 3932 1217 3984
rect 1521 3932 1527 3984
rect 1579 3932 1585 3984
rect 624 3334 630 3386
rect 682 3334 688 3386
rect 1360 3334 1366 3386
rect 1418 3334 1424 3386
rect 49 2736 55 2788
rect 107 2736 113 2788
rect 164 2736 170 2788
rect 222 2736 228 2788
rect 417 2736 423 2788
rect 475 2736 481 2788
rect 785 2736 791 2788
rect 843 2736 849 2788
rect 1153 2736 1159 2788
rect 1211 2736 1217 2788
rect 1521 2736 1527 2788
rect 1579 2736 1585 2788
rect 624 2214 630 2266
rect 682 2214 688 2266
rect 1360 2214 1366 2266
rect 1418 2214 1424 2266
rect 49 1692 55 1744
rect 107 1692 113 1744
rect 164 1692 170 1744
rect 222 1692 228 1744
rect 417 1692 423 1744
rect 475 1692 481 1744
rect 785 1692 791 1744
rect 843 1692 849 1744
rect 1153 1692 1159 1744
rect 1211 1692 1217 1744
rect 1521 1692 1527 1744
rect 1579 1692 1585 1744
rect 624 1094 630 1146
rect 682 1094 688 1146
rect 1360 1094 1366 1146
rect 1418 1094 1424 1146
rect 49 496 55 548
rect 107 496 113 548
rect 164 496 170 548
rect 222 496 228 548
rect 417 496 423 548
rect 475 496 481 548
rect 785 496 791 548
rect 843 496 849 548
rect 1153 496 1159 548
rect 1211 496 1217 548
rect 1521 496 1527 548
rect 1579 496 1585 548
rect 624 -26 630 26
rect 682 -26 688 26
rect 1360 -26 1366 26
rect 1418 -26 1424 26
<< via1 >>
rect 630 10097 682 10106
rect 630 10063 639 10097
rect 639 10063 673 10097
rect 673 10063 682 10097
rect 630 10054 682 10063
rect 1366 10097 1418 10106
rect 1366 10063 1375 10097
rect 1375 10063 1409 10097
rect 1409 10063 1418 10097
rect 1366 10054 1418 10063
rect 55 9499 107 9508
rect 55 9465 64 9499
rect 64 9465 98 9499
rect 98 9465 107 9499
rect 55 9456 107 9465
rect 170 9499 222 9508
rect 170 9465 179 9499
rect 179 9465 213 9499
rect 213 9465 222 9499
rect 170 9456 222 9465
rect 423 9499 475 9508
rect 423 9465 432 9499
rect 432 9465 466 9499
rect 466 9465 475 9499
rect 423 9456 475 9465
rect 791 9499 843 9508
rect 791 9465 800 9499
rect 800 9465 834 9499
rect 834 9465 843 9499
rect 791 9456 843 9465
rect 1159 9499 1211 9508
rect 1159 9465 1168 9499
rect 1168 9465 1202 9499
rect 1202 9465 1211 9499
rect 1159 9456 1211 9465
rect 1527 9499 1579 9508
rect 1527 9465 1536 9499
rect 1536 9465 1570 9499
rect 1570 9465 1579 9499
rect 1527 9456 1579 9465
rect 630 8977 682 8986
rect 630 8943 639 8977
rect 639 8943 673 8977
rect 673 8943 682 8977
rect 630 8934 682 8943
rect 1366 8977 1418 8986
rect 1366 8943 1375 8977
rect 1375 8943 1409 8977
rect 1409 8943 1418 8977
rect 1366 8934 1418 8943
rect 55 8455 107 8464
rect 55 8421 64 8455
rect 64 8421 98 8455
rect 98 8421 107 8455
rect 55 8412 107 8421
rect 170 8455 222 8464
rect 170 8421 179 8455
rect 179 8421 213 8455
rect 213 8421 222 8455
rect 170 8412 222 8421
rect 423 8455 475 8464
rect 423 8421 432 8455
rect 432 8421 466 8455
rect 466 8421 475 8455
rect 423 8412 475 8421
rect 791 8455 843 8464
rect 791 8421 800 8455
rect 800 8421 834 8455
rect 834 8421 843 8455
rect 791 8412 843 8421
rect 1159 8455 1211 8464
rect 1159 8421 1168 8455
rect 1168 8421 1202 8455
rect 1202 8421 1211 8455
rect 1159 8412 1211 8421
rect 1527 8455 1579 8464
rect 1527 8421 1536 8455
rect 1536 8421 1570 8455
rect 1570 8421 1579 8455
rect 1527 8412 1579 8421
rect 630 7857 682 7866
rect 630 7823 639 7857
rect 639 7823 673 7857
rect 673 7823 682 7857
rect 630 7814 682 7823
rect 1366 7857 1418 7866
rect 1366 7823 1375 7857
rect 1375 7823 1409 7857
rect 1409 7823 1418 7857
rect 1366 7814 1418 7823
rect 55 7259 107 7268
rect 55 7225 64 7259
rect 64 7225 98 7259
rect 98 7225 107 7259
rect 55 7216 107 7225
rect 170 7259 222 7268
rect 170 7225 179 7259
rect 179 7225 213 7259
rect 213 7225 222 7259
rect 170 7216 222 7225
rect 423 7259 475 7268
rect 423 7225 432 7259
rect 432 7225 466 7259
rect 466 7225 475 7259
rect 423 7216 475 7225
rect 791 7259 843 7268
rect 791 7225 800 7259
rect 800 7225 834 7259
rect 834 7225 843 7259
rect 791 7216 843 7225
rect 1159 7259 1211 7268
rect 1159 7225 1168 7259
rect 1168 7225 1202 7259
rect 1202 7225 1211 7259
rect 1159 7216 1211 7225
rect 1527 7259 1579 7268
rect 1527 7225 1536 7259
rect 1536 7225 1570 7259
rect 1570 7225 1579 7259
rect 1527 7216 1579 7225
rect 630 6737 682 6746
rect 630 6703 639 6737
rect 639 6703 673 6737
rect 673 6703 682 6737
rect 630 6694 682 6703
rect 1366 6737 1418 6746
rect 1366 6703 1375 6737
rect 1375 6703 1409 6737
rect 1409 6703 1418 6737
rect 1366 6694 1418 6703
rect 55 6215 107 6224
rect 55 6181 64 6215
rect 64 6181 98 6215
rect 98 6181 107 6215
rect 55 6172 107 6181
rect 170 6215 222 6224
rect 170 6181 179 6215
rect 179 6181 213 6215
rect 213 6181 222 6215
rect 170 6172 222 6181
rect 423 6215 475 6224
rect 423 6181 432 6215
rect 432 6181 466 6215
rect 466 6181 475 6215
rect 423 6172 475 6181
rect 791 6215 843 6224
rect 791 6181 800 6215
rect 800 6181 834 6215
rect 834 6181 843 6215
rect 791 6172 843 6181
rect 1159 6215 1211 6224
rect 1159 6181 1168 6215
rect 1168 6181 1202 6215
rect 1202 6181 1211 6215
rect 1159 6172 1211 6181
rect 1527 6215 1579 6224
rect 1527 6181 1536 6215
rect 1536 6181 1570 6215
rect 1570 6181 1579 6215
rect 1527 6172 1579 6181
rect 630 5617 682 5626
rect 630 5583 639 5617
rect 639 5583 673 5617
rect 673 5583 682 5617
rect 630 5574 682 5583
rect 1366 5617 1418 5626
rect 1366 5583 1375 5617
rect 1375 5583 1409 5617
rect 1409 5583 1418 5617
rect 1366 5574 1418 5583
rect 55 5019 107 5028
rect 55 4985 64 5019
rect 64 4985 98 5019
rect 98 4985 107 5019
rect 55 4976 107 4985
rect 170 5019 222 5028
rect 170 4985 179 5019
rect 179 4985 213 5019
rect 213 4985 222 5019
rect 170 4976 222 4985
rect 423 5019 475 5028
rect 423 4985 432 5019
rect 432 4985 466 5019
rect 466 4985 475 5019
rect 423 4976 475 4985
rect 791 5019 843 5028
rect 791 4985 800 5019
rect 800 4985 834 5019
rect 834 4985 843 5019
rect 791 4976 843 4985
rect 1159 5019 1211 5028
rect 1159 4985 1168 5019
rect 1168 4985 1202 5019
rect 1202 4985 1211 5019
rect 1159 4976 1211 4985
rect 1527 5019 1579 5028
rect 1527 4985 1536 5019
rect 1536 4985 1570 5019
rect 1570 4985 1579 5019
rect 1527 4976 1579 4985
rect 630 4497 682 4506
rect 630 4463 639 4497
rect 639 4463 673 4497
rect 673 4463 682 4497
rect 630 4454 682 4463
rect 1366 4497 1418 4506
rect 1366 4463 1375 4497
rect 1375 4463 1409 4497
rect 1409 4463 1418 4497
rect 1366 4454 1418 4463
rect 55 3975 107 3984
rect 55 3941 64 3975
rect 64 3941 98 3975
rect 98 3941 107 3975
rect 55 3932 107 3941
rect 170 3975 222 3984
rect 170 3941 179 3975
rect 179 3941 213 3975
rect 213 3941 222 3975
rect 170 3932 222 3941
rect 423 3975 475 3984
rect 423 3941 432 3975
rect 432 3941 466 3975
rect 466 3941 475 3975
rect 423 3932 475 3941
rect 791 3975 843 3984
rect 791 3941 800 3975
rect 800 3941 834 3975
rect 834 3941 843 3975
rect 791 3932 843 3941
rect 1159 3975 1211 3984
rect 1159 3941 1168 3975
rect 1168 3941 1202 3975
rect 1202 3941 1211 3975
rect 1159 3932 1211 3941
rect 1527 3975 1579 3984
rect 1527 3941 1536 3975
rect 1536 3941 1570 3975
rect 1570 3941 1579 3975
rect 1527 3932 1579 3941
rect 630 3377 682 3386
rect 630 3343 639 3377
rect 639 3343 673 3377
rect 673 3343 682 3377
rect 630 3334 682 3343
rect 1366 3377 1418 3386
rect 1366 3343 1375 3377
rect 1375 3343 1409 3377
rect 1409 3343 1418 3377
rect 1366 3334 1418 3343
rect 55 2779 107 2788
rect 55 2745 64 2779
rect 64 2745 98 2779
rect 98 2745 107 2779
rect 55 2736 107 2745
rect 170 2779 222 2788
rect 170 2745 179 2779
rect 179 2745 213 2779
rect 213 2745 222 2779
rect 170 2736 222 2745
rect 423 2779 475 2788
rect 423 2745 432 2779
rect 432 2745 466 2779
rect 466 2745 475 2779
rect 423 2736 475 2745
rect 791 2779 843 2788
rect 791 2745 800 2779
rect 800 2745 834 2779
rect 834 2745 843 2779
rect 791 2736 843 2745
rect 1159 2779 1211 2788
rect 1159 2745 1168 2779
rect 1168 2745 1202 2779
rect 1202 2745 1211 2779
rect 1159 2736 1211 2745
rect 1527 2779 1579 2788
rect 1527 2745 1536 2779
rect 1536 2745 1570 2779
rect 1570 2745 1579 2779
rect 1527 2736 1579 2745
rect 630 2257 682 2266
rect 630 2223 639 2257
rect 639 2223 673 2257
rect 673 2223 682 2257
rect 630 2214 682 2223
rect 1366 2257 1418 2266
rect 1366 2223 1375 2257
rect 1375 2223 1409 2257
rect 1409 2223 1418 2257
rect 1366 2214 1418 2223
rect 55 1735 107 1744
rect 55 1701 64 1735
rect 64 1701 98 1735
rect 98 1701 107 1735
rect 55 1692 107 1701
rect 170 1735 222 1744
rect 170 1701 179 1735
rect 179 1701 213 1735
rect 213 1701 222 1735
rect 170 1692 222 1701
rect 423 1735 475 1744
rect 423 1701 432 1735
rect 432 1701 466 1735
rect 466 1701 475 1735
rect 423 1692 475 1701
rect 791 1735 843 1744
rect 791 1701 800 1735
rect 800 1701 834 1735
rect 834 1701 843 1735
rect 791 1692 843 1701
rect 1159 1735 1211 1744
rect 1159 1701 1168 1735
rect 1168 1701 1202 1735
rect 1202 1701 1211 1735
rect 1159 1692 1211 1701
rect 1527 1735 1579 1744
rect 1527 1701 1536 1735
rect 1536 1701 1570 1735
rect 1570 1701 1579 1735
rect 1527 1692 1579 1701
rect 630 1137 682 1146
rect 630 1103 639 1137
rect 639 1103 673 1137
rect 673 1103 682 1137
rect 630 1094 682 1103
rect 1366 1137 1418 1146
rect 1366 1103 1375 1137
rect 1375 1103 1409 1137
rect 1409 1103 1418 1137
rect 1366 1094 1418 1103
rect 55 539 107 548
rect 55 505 64 539
rect 64 505 98 539
rect 98 505 107 539
rect 55 496 107 505
rect 170 539 222 548
rect 170 505 179 539
rect 179 505 213 539
rect 213 505 222 539
rect 170 496 222 505
rect 423 539 475 548
rect 423 505 432 539
rect 432 505 466 539
rect 466 505 475 539
rect 423 496 475 505
rect 791 539 843 548
rect 791 505 800 539
rect 800 505 834 539
rect 834 505 843 539
rect 791 496 843 505
rect 1159 539 1211 548
rect 1159 505 1168 539
rect 1168 505 1202 539
rect 1202 505 1211 539
rect 1159 496 1211 505
rect 1527 539 1579 548
rect 1527 505 1536 539
rect 1536 505 1570 539
rect 1570 505 1579 539
rect 1527 496 1579 505
rect 630 17 682 26
rect 630 -17 639 17
rect 639 -17 673 17
rect 673 -17 682 17
rect 630 -26 682 -17
rect 1366 17 1418 26
rect 1366 -17 1375 17
rect 1375 -17 1409 17
rect 1409 -17 1418 17
rect 1366 -26 1418 -17
<< metal2 >>
rect 628 10108 684 10117
rect 628 10043 684 10052
rect 1364 10108 1420 10117
rect 1364 10043 1420 10052
rect 55 9508 107 9514
rect 55 9450 107 9456
rect 168 9510 224 9519
rect 67 8974 95 9450
rect 168 9445 224 9454
rect 421 9510 477 9519
rect 421 9445 477 9454
rect 789 9510 845 9519
rect 789 9445 845 9454
rect 1157 9510 1213 9519
rect 1157 9445 1213 9454
rect 1525 9510 1581 9519
rect 1581 9468 1651 9496
rect 1525 9445 1581 9454
rect 628 8988 684 8997
rect 67 8946 210 8974
rect 182 8475 210 8946
rect 628 8923 684 8932
rect 1364 8988 1420 8997
rect 1364 8923 1420 8932
rect 55 8464 107 8470
rect 55 8406 107 8412
rect 168 8466 224 8475
rect 67 7854 95 8406
rect 168 8401 224 8410
rect 421 8466 477 8475
rect 421 8401 477 8410
rect 789 8466 845 8475
rect 789 8401 845 8410
rect 1157 8466 1213 8475
rect 1157 8401 1213 8410
rect 1525 8466 1581 8475
rect 1525 8401 1581 8410
rect 628 7868 684 7877
rect 67 7826 210 7854
rect 182 7279 210 7826
rect 628 7803 684 7812
rect 1364 7868 1420 7877
rect 1364 7803 1420 7812
rect 55 7268 107 7274
rect 55 7210 107 7216
rect 168 7270 224 7279
rect 67 6734 95 7210
rect 168 7205 224 7214
rect 421 7270 477 7279
rect 421 7205 477 7214
rect 789 7270 845 7279
rect 789 7205 845 7214
rect 1157 7270 1213 7279
rect 1157 7205 1213 7214
rect 1525 7270 1581 7279
rect 1525 7205 1581 7214
rect 628 6748 684 6757
rect 67 6706 210 6734
rect 182 6235 210 6706
rect 628 6683 684 6692
rect 1364 6748 1420 6757
rect 1364 6683 1420 6692
rect 55 6224 107 6230
rect 55 6166 107 6172
rect 168 6226 224 6235
rect 67 5614 95 6166
rect 168 6161 224 6170
rect 421 6226 477 6235
rect 421 6161 477 6170
rect 789 6226 845 6235
rect 789 6161 845 6170
rect 1157 6226 1213 6235
rect 1157 6161 1213 6170
rect 1525 6226 1581 6235
rect 1525 6161 1581 6170
rect 628 5628 684 5637
rect 67 5586 210 5614
rect 182 5039 210 5586
rect 628 5563 684 5572
rect 1364 5628 1420 5637
rect 1364 5563 1420 5572
rect 55 5028 107 5034
rect 55 4970 107 4976
rect 168 5030 224 5039
rect 67 4494 95 4970
rect 168 4965 224 4974
rect 421 5030 477 5039
rect 421 4965 477 4974
rect 789 5030 845 5039
rect 789 4965 845 4974
rect 1157 5030 1213 5039
rect 1157 4965 1213 4974
rect 1525 5030 1581 5039
rect 1525 4965 1581 4974
rect 628 4508 684 4517
rect 67 4466 210 4494
rect 182 3995 210 4466
rect 628 4443 684 4452
rect 1364 4508 1420 4517
rect 1364 4443 1420 4452
rect 55 3984 107 3990
rect 55 3926 107 3932
rect 168 3986 224 3995
rect 67 3374 95 3926
rect 168 3921 224 3930
rect 421 3986 477 3995
rect 421 3921 477 3930
rect 789 3986 845 3995
rect 789 3921 845 3930
rect 1157 3986 1213 3995
rect 1157 3921 1213 3930
rect 1525 3986 1581 3995
rect 1525 3921 1581 3930
rect 628 3388 684 3397
rect 67 3346 210 3374
rect 182 2799 210 3346
rect 628 3323 684 3332
rect 1364 3388 1420 3397
rect 1364 3323 1420 3332
rect 55 2788 107 2794
rect 55 2730 107 2736
rect 168 2790 224 2799
rect 67 2254 95 2730
rect 168 2725 224 2734
rect 421 2790 477 2799
rect 421 2725 477 2734
rect 789 2790 845 2799
rect 789 2725 845 2734
rect 1157 2790 1213 2799
rect 1157 2725 1213 2734
rect 1525 2790 1581 2799
rect 1525 2725 1581 2734
rect 628 2268 684 2277
rect 67 2226 210 2254
rect 182 1755 210 2226
rect 628 2203 684 2212
rect 1364 2268 1420 2277
rect 1364 2203 1420 2212
rect 55 1744 107 1750
rect 55 1686 107 1692
rect 168 1746 224 1755
rect 67 1134 95 1686
rect 168 1681 224 1690
rect 421 1746 477 1755
rect 421 1681 477 1690
rect 789 1746 845 1755
rect 789 1681 845 1690
rect 1157 1746 1213 1755
rect 1157 1681 1213 1690
rect 1525 1746 1581 1755
rect 1525 1681 1581 1690
rect 628 1148 684 1157
rect 67 1106 210 1134
rect 182 559 210 1106
rect 628 1083 684 1092
rect 1364 1148 1420 1157
rect 1364 1083 1420 1092
rect 55 548 107 554
rect 55 490 107 496
rect 168 550 224 559
rect 64 0 92 490
rect 168 485 224 494
rect 421 550 477 559
rect 421 485 477 494
rect 789 550 845 559
rect 789 485 845 494
rect 1157 550 1213 559
rect 1157 485 1213 494
rect 1525 550 1581 559
rect 1525 485 1581 494
rect 628 28 684 37
rect 628 -37 684 -28
rect 1364 28 1420 37
rect 1623 0 1651 9468
rect 1364 -37 1420 -28
<< via2 >>
rect 628 10106 684 10108
rect 628 10054 630 10106
rect 630 10054 682 10106
rect 682 10054 684 10106
rect 628 10052 684 10054
rect 1364 10106 1420 10108
rect 1364 10054 1366 10106
rect 1366 10054 1418 10106
rect 1418 10054 1420 10106
rect 1364 10052 1420 10054
rect 168 9508 224 9510
rect 168 9456 170 9508
rect 170 9456 222 9508
rect 222 9456 224 9508
rect 168 9454 224 9456
rect 421 9508 477 9510
rect 421 9456 423 9508
rect 423 9456 475 9508
rect 475 9456 477 9508
rect 421 9454 477 9456
rect 789 9508 845 9510
rect 789 9456 791 9508
rect 791 9456 843 9508
rect 843 9456 845 9508
rect 789 9454 845 9456
rect 1157 9508 1213 9510
rect 1157 9456 1159 9508
rect 1159 9456 1211 9508
rect 1211 9456 1213 9508
rect 1157 9454 1213 9456
rect 1525 9508 1581 9510
rect 1525 9456 1527 9508
rect 1527 9456 1579 9508
rect 1579 9456 1581 9508
rect 1525 9454 1581 9456
rect 628 8986 684 8988
rect 628 8934 630 8986
rect 630 8934 682 8986
rect 682 8934 684 8986
rect 628 8932 684 8934
rect 1364 8986 1420 8988
rect 1364 8934 1366 8986
rect 1366 8934 1418 8986
rect 1418 8934 1420 8986
rect 1364 8932 1420 8934
rect 168 8464 224 8466
rect 168 8412 170 8464
rect 170 8412 222 8464
rect 222 8412 224 8464
rect 168 8410 224 8412
rect 421 8464 477 8466
rect 421 8412 423 8464
rect 423 8412 475 8464
rect 475 8412 477 8464
rect 421 8410 477 8412
rect 789 8464 845 8466
rect 789 8412 791 8464
rect 791 8412 843 8464
rect 843 8412 845 8464
rect 789 8410 845 8412
rect 1157 8464 1213 8466
rect 1157 8412 1159 8464
rect 1159 8412 1211 8464
rect 1211 8412 1213 8464
rect 1157 8410 1213 8412
rect 1525 8464 1581 8466
rect 1525 8412 1527 8464
rect 1527 8412 1579 8464
rect 1579 8412 1581 8464
rect 1525 8410 1581 8412
rect 628 7866 684 7868
rect 628 7814 630 7866
rect 630 7814 682 7866
rect 682 7814 684 7866
rect 628 7812 684 7814
rect 1364 7866 1420 7868
rect 1364 7814 1366 7866
rect 1366 7814 1418 7866
rect 1418 7814 1420 7866
rect 1364 7812 1420 7814
rect 168 7268 224 7270
rect 168 7216 170 7268
rect 170 7216 222 7268
rect 222 7216 224 7268
rect 168 7214 224 7216
rect 421 7268 477 7270
rect 421 7216 423 7268
rect 423 7216 475 7268
rect 475 7216 477 7268
rect 421 7214 477 7216
rect 789 7268 845 7270
rect 789 7216 791 7268
rect 791 7216 843 7268
rect 843 7216 845 7268
rect 789 7214 845 7216
rect 1157 7268 1213 7270
rect 1157 7216 1159 7268
rect 1159 7216 1211 7268
rect 1211 7216 1213 7268
rect 1157 7214 1213 7216
rect 1525 7268 1581 7270
rect 1525 7216 1527 7268
rect 1527 7216 1579 7268
rect 1579 7216 1581 7268
rect 1525 7214 1581 7216
rect 628 6746 684 6748
rect 628 6694 630 6746
rect 630 6694 682 6746
rect 682 6694 684 6746
rect 628 6692 684 6694
rect 1364 6746 1420 6748
rect 1364 6694 1366 6746
rect 1366 6694 1418 6746
rect 1418 6694 1420 6746
rect 1364 6692 1420 6694
rect 168 6224 224 6226
rect 168 6172 170 6224
rect 170 6172 222 6224
rect 222 6172 224 6224
rect 168 6170 224 6172
rect 421 6224 477 6226
rect 421 6172 423 6224
rect 423 6172 475 6224
rect 475 6172 477 6224
rect 421 6170 477 6172
rect 789 6224 845 6226
rect 789 6172 791 6224
rect 791 6172 843 6224
rect 843 6172 845 6224
rect 789 6170 845 6172
rect 1157 6224 1213 6226
rect 1157 6172 1159 6224
rect 1159 6172 1211 6224
rect 1211 6172 1213 6224
rect 1157 6170 1213 6172
rect 1525 6224 1581 6226
rect 1525 6172 1527 6224
rect 1527 6172 1579 6224
rect 1579 6172 1581 6224
rect 1525 6170 1581 6172
rect 628 5626 684 5628
rect 628 5574 630 5626
rect 630 5574 682 5626
rect 682 5574 684 5626
rect 628 5572 684 5574
rect 1364 5626 1420 5628
rect 1364 5574 1366 5626
rect 1366 5574 1418 5626
rect 1418 5574 1420 5626
rect 1364 5572 1420 5574
rect 168 5028 224 5030
rect 168 4976 170 5028
rect 170 4976 222 5028
rect 222 4976 224 5028
rect 168 4974 224 4976
rect 421 5028 477 5030
rect 421 4976 423 5028
rect 423 4976 475 5028
rect 475 4976 477 5028
rect 421 4974 477 4976
rect 789 5028 845 5030
rect 789 4976 791 5028
rect 791 4976 843 5028
rect 843 4976 845 5028
rect 789 4974 845 4976
rect 1157 5028 1213 5030
rect 1157 4976 1159 5028
rect 1159 4976 1211 5028
rect 1211 4976 1213 5028
rect 1157 4974 1213 4976
rect 1525 5028 1581 5030
rect 1525 4976 1527 5028
rect 1527 4976 1579 5028
rect 1579 4976 1581 5028
rect 1525 4974 1581 4976
rect 628 4506 684 4508
rect 628 4454 630 4506
rect 630 4454 682 4506
rect 682 4454 684 4506
rect 628 4452 684 4454
rect 1364 4506 1420 4508
rect 1364 4454 1366 4506
rect 1366 4454 1418 4506
rect 1418 4454 1420 4506
rect 1364 4452 1420 4454
rect 168 3984 224 3986
rect 168 3932 170 3984
rect 170 3932 222 3984
rect 222 3932 224 3984
rect 168 3930 224 3932
rect 421 3984 477 3986
rect 421 3932 423 3984
rect 423 3932 475 3984
rect 475 3932 477 3984
rect 421 3930 477 3932
rect 789 3984 845 3986
rect 789 3932 791 3984
rect 791 3932 843 3984
rect 843 3932 845 3984
rect 789 3930 845 3932
rect 1157 3984 1213 3986
rect 1157 3932 1159 3984
rect 1159 3932 1211 3984
rect 1211 3932 1213 3984
rect 1157 3930 1213 3932
rect 1525 3984 1581 3986
rect 1525 3932 1527 3984
rect 1527 3932 1579 3984
rect 1579 3932 1581 3984
rect 1525 3930 1581 3932
rect 628 3386 684 3388
rect 628 3334 630 3386
rect 630 3334 682 3386
rect 682 3334 684 3386
rect 628 3332 684 3334
rect 1364 3386 1420 3388
rect 1364 3334 1366 3386
rect 1366 3334 1418 3386
rect 1418 3334 1420 3386
rect 1364 3332 1420 3334
rect 168 2788 224 2790
rect 168 2736 170 2788
rect 170 2736 222 2788
rect 222 2736 224 2788
rect 168 2734 224 2736
rect 421 2788 477 2790
rect 421 2736 423 2788
rect 423 2736 475 2788
rect 475 2736 477 2788
rect 421 2734 477 2736
rect 789 2788 845 2790
rect 789 2736 791 2788
rect 791 2736 843 2788
rect 843 2736 845 2788
rect 789 2734 845 2736
rect 1157 2788 1213 2790
rect 1157 2736 1159 2788
rect 1159 2736 1211 2788
rect 1211 2736 1213 2788
rect 1157 2734 1213 2736
rect 1525 2788 1581 2790
rect 1525 2736 1527 2788
rect 1527 2736 1579 2788
rect 1579 2736 1581 2788
rect 1525 2734 1581 2736
rect 628 2266 684 2268
rect 628 2214 630 2266
rect 630 2214 682 2266
rect 682 2214 684 2266
rect 628 2212 684 2214
rect 1364 2266 1420 2268
rect 1364 2214 1366 2266
rect 1366 2214 1418 2266
rect 1418 2214 1420 2266
rect 1364 2212 1420 2214
rect 168 1744 224 1746
rect 168 1692 170 1744
rect 170 1692 222 1744
rect 222 1692 224 1744
rect 168 1690 224 1692
rect 421 1744 477 1746
rect 421 1692 423 1744
rect 423 1692 475 1744
rect 475 1692 477 1744
rect 421 1690 477 1692
rect 789 1744 845 1746
rect 789 1692 791 1744
rect 791 1692 843 1744
rect 843 1692 845 1744
rect 789 1690 845 1692
rect 1157 1744 1213 1746
rect 1157 1692 1159 1744
rect 1159 1692 1211 1744
rect 1211 1692 1213 1744
rect 1157 1690 1213 1692
rect 1525 1744 1581 1746
rect 1525 1692 1527 1744
rect 1527 1692 1579 1744
rect 1579 1692 1581 1744
rect 1525 1690 1581 1692
rect 628 1146 684 1148
rect 628 1094 630 1146
rect 630 1094 682 1146
rect 682 1094 684 1146
rect 628 1092 684 1094
rect 1364 1146 1420 1148
rect 1364 1094 1366 1146
rect 1366 1094 1418 1146
rect 1418 1094 1420 1146
rect 1364 1092 1420 1094
rect 168 548 224 550
rect 168 496 170 548
rect 170 496 222 548
rect 222 496 224 548
rect 168 494 224 496
rect 421 548 477 550
rect 421 496 423 548
rect 423 496 475 548
rect 475 496 477 548
rect 421 494 477 496
rect 789 548 845 550
rect 789 496 791 548
rect 791 496 843 548
rect 843 496 845 548
rect 789 494 845 496
rect 1157 548 1213 550
rect 1157 496 1159 548
rect 1159 496 1211 548
rect 1211 496 1213 548
rect 1157 494 1213 496
rect 1525 548 1581 550
rect 1525 496 1527 548
rect 1527 496 1579 548
rect 1579 496 1581 548
rect 1525 494 1581 496
rect 628 26 684 28
rect 628 -26 630 26
rect 630 -26 682 26
rect 682 -26 684 26
rect 628 -28 684 -26
rect 1364 26 1420 28
rect 1364 -26 1366 26
rect 1366 -26 1418 26
rect 1418 -26 1420 26
rect 1364 -28 1420 -26
<< metal3 >>
rect 607 10108 705 10129
rect 607 10052 628 10108
rect 684 10052 705 10108
rect 607 10031 705 10052
rect 1343 10108 1441 10129
rect 1343 10052 1364 10108
rect 1420 10052 1441 10108
rect 1343 10031 1441 10052
rect 163 9512 229 9515
rect 416 9512 482 9515
rect 784 9512 850 9515
rect 1152 9512 1218 9515
rect 1520 9512 1586 9515
rect 163 9510 1586 9512
rect 163 9454 168 9510
rect 224 9454 421 9510
rect 477 9454 789 9510
rect 845 9454 1157 9510
rect 1213 9454 1525 9510
rect 1581 9454 1586 9510
rect 163 9452 1586 9454
rect 163 9449 229 9452
rect 416 9449 482 9452
rect 784 9449 850 9452
rect 1152 9449 1218 9452
rect 1520 9449 1586 9452
rect 607 8988 705 9009
rect 607 8932 628 8988
rect 684 8932 705 8988
rect 607 8911 705 8932
rect 1343 8988 1441 9009
rect 1343 8932 1364 8988
rect 1420 8932 1441 8988
rect 1343 8911 1441 8932
rect 163 8468 229 8471
rect 416 8468 482 8471
rect 784 8468 850 8471
rect 1152 8468 1218 8471
rect 1520 8468 1586 8471
rect 163 8466 1586 8468
rect 163 8410 168 8466
rect 224 8410 421 8466
rect 477 8410 789 8466
rect 845 8410 1157 8466
rect 1213 8410 1525 8466
rect 1581 8410 1586 8466
rect 163 8408 1586 8410
rect 163 8405 229 8408
rect 416 8405 482 8408
rect 784 8405 850 8408
rect 1152 8405 1218 8408
rect 1520 8405 1586 8408
rect 607 7868 705 7889
rect 607 7812 628 7868
rect 684 7812 705 7868
rect 607 7791 705 7812
rect 1343 7868 1441 7889
rect 1343 7812 1364 7868
rect 1420 7812 1441 7868
rect 1343 7791 1441 7812
rect 163 7272 229 7275
rect 416 7272 482 7275
rect 784 7272 850 7275
rect 1152 7272 1218 7275
rect 1520 7272 1586 7275
rect 163 7270 1586 7272
rect 163 7214 168 7270
rect 224 7214 421 7270
rect 477 7214 789 7270
rect 845 7214 1157 7270
rect 1213 7214 1525 7270
rect 1581 7214 1586 7270
rect 163 7212 1586 7214
rect 163 7209 229 7212
rect 416 7209 482 7212
rect 784 7209 850 7212
rect 1152 7209 1218 7212
rect 1520 7209 1586 7212
rect 607 6748 705 6769
rect 607 6692 628 6748
rect 684 6692 705 6748
rect 607 6671 705 6692
rect 1343 6748 1441 6769
rect 1343 6692 1364 6748
rect 1420 6692 1441 6748
rect 1343 6671 1441 6692
rect 163 6228 229 6231
rect 416 6228 482 6231
rect 784 6228 850 6231
rect 1152 6228 1218 6231
rect 1520 6228 1586 6231
rect 163 6226 1586 6228
rect 163 6170 168 6226
rect 224 6170 421 6226
rect 477 6170 789 6226
rect 845 6170 1157 6226
rect 1213 6170 1525 6226
rect 1581 6170 1586 6226
rect 163 6168 1586 6170
rect 163 6165 229 6168
rect 416 6165 482 6168
rect 784 6165 850 6168
rect 1152 6165 1218 6168
rect 1520 6165 1586 6168
rect 607 5628 705 5649
rect 607 5572 628 5628
rect 684 5572 705 5628
rect 607 5551 705 5572
rect 1343 5628 1441 5649
rect 1343 5572 1364 5628
rect 1420 5572 1441 5628
rect 1343 5551 1441 5572
rect 163 5032 229 5035
rect 416 5032 482 5035
rect 784 5032 850 5035
rect 1152 5032 1218 5035
rect 1520 5032 1586 5035
rect 163 5030 1586 5032
rect 163 4974 168 5030
rect 224 4974 421 5030
rect 477 4974 789 5030
rect 845 4974 1157 5030
rect 1213 4974 1525 5030
rect 1581 4974 1586 5030
rect 163 4972 1586 4974
rect 163 4969 229 4972
rect 416 4969 482 4972
rect 784 4969 850 4972
rect 1152 4969 1218 4972
rect 1520 4969 1586 4972
rect 607 4508 705 4529
rect 607 4452 628 4508
rect 684 4452 705 4508
rect 607 4431 705 4452
rect 1343 4508 1441 4529
rect 1343 4452 1364 4508
rect 1420 4452 1441 4508
rect 1343 4431 1441 4452
rect 163 3988 229 3991
rect 416 3988 482 3991
rect 784 3988 850 3991
rect 1152 3988 1218 3991
rect 1520 3988 1586 3991
rect 163 3986 1586 3988
rect 163 3930 168 3986
rect 224 3930 421 3986
rect 477 3930 789 3986
rect 845 3930 1157 3986
rect 1213 3930 1525 3986
rect 1581 3930 1586 3986
rect 163 3928 1586 3930
rect 163 3925 229 3928
rect 416 3925 482 3928
rect 784 3925 850 3928
rect 1152 3925 1218 3928
rect 1520 3925 1586 3928
rect 607 3388 705 3409
rect 607 3332 628 3388
rect 684 3332 705 3388
rect 607 3311 705 3332
rect 1343 3388 1441 3409
rect 1343 3332 1364 3388
rect 1420 3332 1441 3388
rect 1343 3311 1441 3332
rect 163 2792 229 2795
rect 416 2792 482 2795
rect 784 2792 850 2795
rect 1152 2792 1218 2795
rect 1520 2792 1586 2795
rect 163 2790 1586 2792
rect 163 2734 168 2790
rect 224 2734 421 2790
rect 477 2734 789 2790
rect 845 2734 1157 2790
rect 1213 2734 1525 2790
rect 1581 2734 1586 2790
rect 163 2732 1586 2734
rect 163 2729 229 2732
rect 416 2729 482 2732
rect 784 2729 850 2732
rect 1152 2729 1218 2732
rect 1520 2729 1586 2732
rect 607 2268 705 2289
rect 607 2212 628 2268
rect 684 2212 705 2268
rect 607 2191 705 2212
rect 1343 2268 1441 2289
rect 1343 2212 1364 2268
rect 1420 2212 1441 2268
rect 1343 2191 1441 2212
rect 163 1748 229 1751
rect 416 1748 482 1751
rect 784 1748 850 1751
rect 1152 1748 1218 1751
rect 1520 1748 1586 1751
rect 163 1746 1586 1748
rect 163 1690 168 1746
rect 224 1690 421 1746
rect 477 1690 789 1746
rect 845 1690 1157 1746
rect 1213 1690 1525 1746
rect 1581 1690 1586 1746
rect 163 1688 1586 1690
rect 163 1685 229 1688
rect 416 1685 482 1688
rect 784 1685 850 1688
rect 1152 1685 1218 1688
rect 1520 1685 1586 1688
rect 607 1148 705 1169
rect 607 1092 628 1148
rect 684 1092 705 1148
rect 607 1071 705 1092
rect 1343 1148 1441 1169
rect 1343 1092 1364 1148
rect 1420 1092 1441 1148
rect 1343 1071 1441 1092
rect 163 552 229 555
rect 416 552 482 555
rect 784 552 850 555
rect 1152 552 1218 555
rect 1520 552 1586 555
rect 163 550 1586 552
rect 163 494 168 550
rect 224 494 421 550
rect 477 494 789 550
rect 845 494 1157 550
rect 1213 494 1525 550
rect 1581 494 1586 550
rect 163 492 1586 494
rect 163 489 229 492
rect 416 489 482 492
rect 784 489 850 492
rect 1152 489 1218 492
rect 1520 489 1586 492
rect 607 28 705 49
rect 607 -28 628 28
rect 684 -28 705 28
rect 607 -49 705 -28
rect 1343 28 1441 49
rect 1343 -28 1364 28
rect 1420 -28 1441 28
rect 1343 -49 1441 -28
use contact_9  contact_9_18
timestamp 1636140361
transform 1 0 163 0 1 485
box 0 0 1 1
use contact_8  contact_8_20
timestamp 1636140361
transform 1 0 49 0 1 490
box 0 0 1 1
use contact_7  contact_7_20
timestamp 1636140361
transform 1 0 52 0 1 489
box 0 0 1 1
use contact_8  contact_8_21
timestamp 1636140361
transform 1 0 164 0 1 490
box 0 0 1 1
use contact_7  contact_7_21
timestamp 1636140361
transform 1 0 167 0 1 489
box 0 0 1 1
use contact_8  contact_8_22
timestamp 1636140361
transform 1 0 49 0 1 490
box 0 0 1 1
use contact_7  contact_7_22
timestamp 1636140361
transform 1 0 52 0 1 489
box 0 0 1 1
use pinv_20  pinv_20_4
timestamp 1636140361
transform 1 0 368 0 -1 2240
box -36 -17 404 1177
use pinv_20  pinv_20_5
timestamp 1636140361
transform 1 0 0 0 -1 2240
box -36 -17 404 1177
use pinv_20  pinv_20_6
timestamp 1636140361
transform 1 0 368 0 1 0
box -36 -17 404 1177
use pinv_20  pinv_20_7
timestamp 1636140361
transform 1 0 0 0 1 0
box -36 -17 404 1177
use contact_8  contact_8_9
timestamp 1636140361
transform 1 0 785 0 1 490
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1636140361
transform 1 0 788 0 1 489
box 0 0 1 1
use contact_9  contact_9_10
timestamp 1636140361
transform 1 0 416 0 1 485
box 0 0 1 1
use contact_8  contact_8_11
timestamp 1636140361
transform 1 0 417 0 1 490
box 0 0 1 1
use contact_7  contact_7_11
timestamp 1636140361
transform 1 0 420 0 1 489
box 0 0 1 1
use contact_9  contact_9_11
timestamp 1636140361
transform 1 0 623 0 1 -37
box 0 0 1 1
use contact_8  contact_8_13
timestamp 1636140361
transform 1 0 624 0 1 -32
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1636140361
transform 1 0 627 0 1 -33
box 0 0 1 1
use contact_9  contact_9_19
timestamp 1636140361
transform 1 0 784 0 1 485
box 0 0 1 1
use contact_9  contact_9_9
timestamp 1636140361
transform 1 0 623 0 1 1083
box 0 0 1 1
use contact_8  contact_8_12
timestamp 1636140361
transform 1 0 624 0 1 1088
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1636140361
transform 1 0 627 0 1 1087
box 0 0 1 1
use contact_9  contact_9_12
timestamp 1636140361
transform 1 0 623 0 1 1083
box 0 0 1 1
use contact_8  contact_8_14
timestamp 1636140361
transform 1 0 624 0 1 1088
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1636140361
transform 1 0 627 0 1 1087
box 0 0 1 1
use pinv_20  pinv_20_16
timestamp 1636140361
transform 1 0 736 0 1 0
box -36 -17 404 1177
use pinv_20  pinv_20_19
timestamp 1636140361
transform 1 0 736 0 -1 2240
box -36 -17 404 1177
use contact_9  contact_9_7
timestamp 1636140361
transform 1 0 1152 0 1 485
box 0 0 1 1
use pinv_20  pinv_20_3
timestamp 1636140361
transform 1 0 1104 0 -1 2240
box -36 -17 404 1177
use pinv_20  pinv_20_0
timestamp 1636140361
transform 1 0 1104 0 1 0
box -36 -17 404 1177
use contact_7  contact_7_1
timestamp 1636140361
transform 1 0 1156 0 1 489
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1636140361
transform 1 0 1153 0 1 490
box 0 0 1 1
use contact_9  contact_9_0
timestamp 1636140361
transform 1 0 1520 0 1 485
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1636140361
transform 1 0 1359 0 1 -37
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1636140361
transform 1 0 1360 0 1 -32
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1636140361
transform 1 0 1363 0 1 -33
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1636140361
transform 1 0 1521 0 1 490
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1636140361
transform 1 0 1524 0 1 489
box 0 0 1 1
use contact_7  contact_7_0
timestamp 1636140361
transform 1 0 1363 0 1 1087
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1636140361
transform 1 0 1359 0 1 1083
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1636140361
transform 1 0 1360 0 1 1088
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1636140361
transform 1 0 1363 0 1 1087
box 0 0 1 1
use contact_9  contact_9_8
timestamp 1636140361
transform 1 0 1359 0 1 1083
box 0 0 1 1
use contact_8  contact_8_8
timestamp 1636140361
transform 1 0 1360 0 1 1088
box 0 0 1 1
use pinv_20  pinv_20_1
timestamp 1636140361
transform 1 0 1472 0 1 0
box -36 -17 404 1177
use pinv_20  pinv_20_2
timestamp 1636140361
transform 1 0 1472 0 -1 2240
box -36 -17 404 1177
use pinv_20  pinv_20_15
timestamp 1636140361
transform 1 0 0 0 1 2240
box -36 -17 404 1177
use pinv_20  pinv_20_14
timestamp 1636140361
transform 1 0 368 0 1 2240
box -36 -17 404 1177
use contact_7  contact_7_17
timestamp 1636140361
transform 1 0 52 0 1 1685
box 0 0 1 1
use contact_8  contact_8_17
timestamp 1636140361
transform 1 0 49 0 1 1686
box 0 0 1 1
use contact_7  contact_7_16
timestamp 1636140361
transform 1 0 167 0 1 1685
box 0 0 1 1
use contact_8  contact_8_16
timestamp 1636140361
transform 1 0 164 0 1 1686
box 0 0 1 1
use contact_9  contact_9_15
timestamp 1636140361
transform 1 0 163 0 1 1681
box 0 0 1 1
use contact_9  contact_9_16
timestamp 1636140361
transform 1 0 784 0 1 1681
box 0 0 1 1
use contact_8  contact_8_18
timestamp 1636140361
transform 1 0 785 0 1 1686
box 0 0 1 1
use contact_7  contact_7_18
timestamp 1636140361
transform 1 0 788 0 1 1685
box 0 0 1 1
use contact_9  contact_9_17
timestamp 1636140361
transform 1 0 416 0 1 1681
box 0 0 1 1
use contact_8  contact_8_19
timestamp 1636140361
transform 1 0 417 0 1 1686
box 0 0 1 1
use contact_7  contact_7_19
timestamp 1636140361
transform 1 0 420 0 1 1685
box 0 0 1 1
use contact_8  contact_8_10
timestamp 1636140361
transform 1 0 624 0 1 2208
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1636140361
transform 1 0 627 0 1 2207
box 0 0 1 1
use contact_9  contact_9_13
timestamp 1636140361
transform 1 0 623 0 1 2203
box 0 0 1 1
use contact_8  contact_8_15
timestamp 1636140361
transform 1 0 624 0 1 2208
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1636140361
transform 1 0 627 0 1 2207
box 0 0 1 1
use contact_9  contact_9_14
timestamp 1636140361
transform 1 0 623 0 1 2203
box 0 0 1 1
use pinv_20  pinv_20_18
timestamp 1636140361
transform 1 0 736 0 1 2240
box -36 -17 404 1177
use pinv_20  pinv_20_13
timestamp 1636140361
transform 1 0 1104 0 1 2240
box -36 -17 404 1177
use contact_7  contact_7_8
timestamp 1636140361
transform 1 0 1156 0 1 1685
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1636140361
transform 1 0 1153 0 1 1686
box 0 0 1 1
use contact_9  contact_9_5
timestamp 1636140361
transform 1 0 1152 0 1 1681
box 0 0 1 1
use contact_9  contact_9_4
timestamp 1636140361
transform 1 0 1520 0 1 1681
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1636140361
transform 1 0 1521 0 1 1686
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1636140361
transform 1 0 1524 0 1 1685
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1636140361
transform 1 0 1359 0 1 2203
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1636140361
transform 1 0 1360 0 1 2208
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1636140361
transform 1 0 1363 0 1 2207
box 0 0 1 1
use contact_9  contact_9_6
timestamp 1636140361
transform 1 0 1359 0 1 2203
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1636140361
transform 1 0 1360 0 1 2208
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1636140361
transform 1 0 1363 0 1 2207
box 0 0 1 1
use pinv_20  pinv_20_12
timestamp 1636140361
transform 1 0 1472 0 1 2240
box -36 -17 404 1177
use pinv_20  pinv_20_9
timestamp 1636140361
transform 1 0 0 0 -1 4480
box -36 -17 404 1177
use pinv_20  pinv_20_8
timestamp 1636140361
transform 1 0 368 0 -1 4480
box -36 -17 404 1177
use contact_7  contact_7_27
timestamp 1636140361
transform 1 0 52 0 1 2729
box 0 0 1 1
use contact_8  contact_8_26
timestamp 1636140361
transform 1 0 49 0 1 2730
box 0 0 1 1
use contact_7  contact_7_26
timestamp 1636140361
transform 1 0 167 0 1 2729
box 0 0 1 1
use contact_8  contact_8_25
timestamp 1636140361
transform 1 0 164 0 1 2730
box 0 0 1 1
use contact_9  contact_9_22
timestamp 1636140361
transform 1 0 163 0 1 2725
box 0 0 1 1
use contact_9  contact_9_23
timestamp 1636140361
transform 1 0 784 0 1 2725
box 0 0 1 1
use contact_8  contact_8_27
timestamp 1636140361
transform 1 0 785 0 1 2730
box 0 0 1 1
use contact_7  contact_7_28
timestamp 1636140361
transform 1 0 788 0 1 2729
box 0 0 1 1
use contact_9  contact_9_24
timestamp 1636140361
transform 1 0 416 0 1 2725
box 0 0 1 1
use contact_8  contact_8_28
timestamp 1636140361
transform 1 0 417 0 1 2730
box 0 0 1 1
use contact_7  contact_7_29
timestamp 1636140361
transform 1 0 420 0 1 2729
box 0 0 1 1
use contact_9  contact_9_27
timestamp 1636140361
transform 1 0 623 0 1 3323
box 0 0 1 1
use contact_8  contact_8_31
timestamp 1636140361
transform 1 0 624 0 1 3328
box 0 0 1 1
use contact_7  contact_7_32
timestamp 1636140361
transform 1 0 627 0 1 3327
box 0 0 1 1
use contact_9  contact_9_28
timestamp 1636140361
transform 1 0 623 0 1 3323
box 0 0 1 1
use contact_8  contact_8_32
timestamp 1636140361
transform 1 0 624 0 1 3328
box 0 0 1 1
use contact_7  contact_7_33
timestamp 1636140361
transform 1 0 627 0 1 3327
box 0 0 1 1
use pinv_20  pinv_20_17
timestamp 1636140361
transform 1 0 736 0 -1 4480
box -36 -17 404 1177
use pinv_20  pinv_20_10
timestamp 1636140361
transform 1 0 1104 0 -1 4480
box -36 -17 404 1177
use contact_7  contact_7_47
timestamp 1636140361
transform 1 0 1156 0 1 2729
box 0 0 1 1
use contact_8  contact_8_47
timestamp 1636140361
transform 1 0 1153 0 1 2730
box 0 0 1 1
use contact_9  contact_9_38
timestamp 1636140361
transform 1 0 1152 0 1 2725
box 0 0 1 1
use contact_9  contact_9_37
timestamp 1636140361
transform 1 0 1520 0 1 2725
box 0 0 1 1
use contact_8  contact_8_44
timestamp 1636140361
transform 1 0 1521 0 1 2730
box 0 0 1 1
use contact_7  contact_7_44
timestamp 1636140361
transform 1 0 1524 0 1 2729
box 0 0 1 1
use contact_9  contact_9_34
timestamp 1636140361
transform 1 0 1359 0 1 3323
box 0 0 1 1
use contact_8  contact_8_41
timestamp 1636140361
transform 1 0 1360 0 1 3328
box 0 0 1 1
use contact_7  contact_7_41
timestamp 1636140361
transform 1 0 1363 0 1 3327
box 0 0 1 1
use contact_9  contact_9_36
timestamp 1636140361
transform 1 0 1359 0 1 3323
box 0 0 1 1
use contact_8  contact_8_43
timestamp 1636140361
transform 1 0 1360 0 1 3328
box 0 0 1 1
use contact_7  contact_7_43
timestamp 1636140361
transform 1 0 1363 0 1 3327
box 0 0 1 1
use pinv_20  pinv_20_11
timestamp 1636140361
transform 1 0 1472 0 -1 4480
box -36 -17 404 1177
use pinv_20  pinv_20_44
timestamp 1636140361
transform 1 0 0 0 1 4480
box -36 -17 404 1177
use pinv_20  pinv_20_43
timestamp 1636140361
transform 1 0 368 0 1 4480
box -36 -17 404 1177
use contact_8  contact_8_38
timestamp 1636140361
transform 1 0 49 0 1 3926
box 0 0 1 1
use contact_7  contact_7_38
timestamp 1636140361
transform 1 0 167 0 1 3925
box 0 0 1 1
use contact_8  contact_8_37
timestamp 1636140361
transform 1 0 164 0 1 3926
box 0 0 1 1
use contact_9  contact_9_32
timestamp 1636140361
transform 1 0 163 0 1 3921
box 0 0 1 1
use contact_7  contact_7_23
timestamp 1636140361
transform 1 0 52 0 1 3925
box 0 0 1 1
use contact_9  contact_9_20
timestamp 1636140361
transform 1 0 784 0 1 3921
box 0 0 1 1
use contact_8  contact_8_23
timestamp 1636140361
transform 1 0 785 0 1 3926
box 0 0 1 1
use contact_7  contact_7_24
timestamp 1636140361
transform 1 0 788 0 1 3925
box 0 0 1 1
use contact_9  contact_9_21
timestamp 1636140361
transform 1 0 416 0 1 3921
box 0 0 1 1
use contact_8  contact_8_24
timestamp 1636140361
transform 1 0 417 0 1 3926
box 0 0 1 1
use contact_7  contact_7_25
timestamp 1636140361
transform 1 0 420 0 1 3925
box 0 0 1 1
use contact_9  contact_9_25
timestamp 1636140361
transform 1 0 623 0 1 4443
box 0 0 1 1
use contact_8  contact_8_29
timestamp 1636140361
transform 1 0 624 0 1 4448
box 0 0 1 1
use contact_7  contact_7_30
timestamp 1636140361
transform 1 0 627 0 1 4447
box 0 0 1 1
use contact_9  contact_9_26
timestamp 1636140361
transform 1 0 623 0 1 4443
box 0 0 1 1
use contact_8  contact_8_30
timestamp 1636140361
transform 1 0 624 0 1 4448
box 0 0 1 1
use contact_7  contact_7_31
timestamp 1636140361
transform 1 0 627 0 1 4447
box 0 0 1 1
use pinv_20  pinv_20_42
timestamp 1636140361
transform 1 0 736 0 1 4480
box -36 -17 404 1177
use pinv_20  pinv_20_41
timestamp 1636140361
transform 1 0 1104 0 1 4480
box -36 -17 404 1177
use contact_7  contact_7_42
timestamp 1636140361
transform 1 0 1156 0 1 3925
box 0 0 1 1
use contact_8  contact_8_42
timestamp 1636140361
transform 1 0 1153 0 1 3926
box 0 0 1 1
use contact_9  contact_9_35
timestamp 1636140361
transform 1 0 1152 0 1 3921
box 0 0 1 1
use contact_9  contact_9_33
timestamp 1636140361
transform 1 0 1520 0 1 3921
box 0 0 1 1
use contact_8  contact_8_40
timestamp 1636140361
transform 1 0 1521 0 1 3926
box 0 0 1 1
use contact_7  contact_7_40
timestamp 1636140361
transform 1 0 1524 0 1 3925
box 0 0 1 1
use contact_8  contact_8_39
timestamp 1636140361
transform 1 0 1360 0 1 4448
box 0 0 1 1
use contact_7  contact_7_39
timestamp 1636140361
transform 1 0 1363 0 1 4447
box 0 0 1 1
use contact_9  contact_9_41
timestamp 1636140361
transform 1 0 1359 0 1 4443
box 0 0 1 1
use contact_8  contact_8_48
timestamp 1636140361
transform 1 0 1360 0 1 4448
box 0 0 1 1
use contact_7  contact_7_48
timestamp 1636140361
transform 1 0 1363 0 1 4447
box 0 0 1 1
use contact_9  contact_9_42
timestamp 1636140361
transform 1 0 1359 0 1 4443
box 0 0 1 1
use pinv_20  pinv_20_40
timestamp 1636140361
transform 1 0 1472 0 1 4480
box -36 -17 404 1177
use pinv_20  pinv_20_23
timestamp 1636140361
transform 1 0 368 0 -1 6720
box -36 -17 404 1177
use pinv_20  pinv_20_22
timestamp 1636140361
transform 1 0 0 0 -1 6720
box -36 -17 404 1177
use contact_7  contact_7_35
timestamp 1636140361
transform 1 0 52 0 1 4969
box 0 0 1 1
use contact_8  contact_8_34
timestamp 1636140361
transform 1 0 49 0 1 4970
box 0 0 1 1
use contact_7  contact_7_34
timestamp 1636140361
transform 1 0 167 0 1 4969
box 0 0 1 1
use contact_8  contact_8_33
timestamp 1636140361
transform 1 0 164 0 1 4970
box 0 0 1 1
use contact_9  contact_9_29
timestamp 1636140361
transform 1 0 163 0 1 4965
box 0 0 1 1
use contact_9  contact_9_30
timestamp 1636140361
transform 1 0 784 0 1 4965
box 0 0 1 1
use contact_8  contact_8_35
timestamp 1636140361
transform 1 0 785 0 1 4970
box 0 0 1 1
use contact_7  contact_7_36
timestamp 1636140361
transform 1 0 788 0 1 4969
box 0 0 1 1
use contact_9  contact_9_31
timestamp 1636140361
transform 1 0 416 0 1 4965
box 0 0 1 1
use contact_8  contact_8_36
timestamp 1636140361
transform 1 0 417 0 1 4970
box 0 0 1 1
use contact_7  contact_7_37
timestamp 1636140361
transform 1 0 420 0 1 4969
box 0 0 1 1
use contact_9  contact_9_55
timestamp 1636140361
transform 1 0 623 0 1 5563
box 0 0 1 1
use contact_8  contact_8_62
timestamp 1636140361
transform 1 0 624 0 1 5568
box 0 0 1 1
use contact_7  contact_7_61
timestamp 1636140361
transform 1 0 627 0 1 5567
box 0 0 1 1
use contact_9  contact_9_58
timestamp 1636140361
transform 1 0 623 0 1 5563
box 0 0 1 1
use contact_8  contact_8_65
timestamp 1636140361
transform 1 0 624 0 1 5568
box 0 0 1 1
use contact_7  contact_7_68
timestamp 1636140361
transform 1 0 627 0 1 5567
box 0 0 1 1
use pinv_20  pinv_20_39
timestamp 1636140361
transform 1 0 736 0 -1 6720
box -36 -17 404 1177
use pinv_20  pinv_20_20
timestamp 1636140361
transform 1 0 1104 0 -1 6720
box -36 -17 404 1177
use contact_7  contact_7_46
timestamp 1636140361
transform 1 0 1156 0 1 4969
box 0 0 1 1
use contact_8  contact_8_46
timestamp 1636140361
transform 1 0 1153 0 1 4970
box 0 0 1 1
use contact_9  contact_9_40
timestamp 1636140361
transform 1 0 1152 0 1 4965
box 0 0 1 1
use contact_9  contact_9_39
timestamp 1636140361
transform 1 0 1520 0 1 4965
box 0 0 1 1
use contact_8  contact_8_45
timestamp 1636140361
transform 1 0 1521 0 1 4970
box 0 0 1 1
use contact_7  contact_7_45
timestamp 1636140361
transform 1 0 1524 0 1 4969
box 0 0 1 1
use contact_7  contact_7_49
timestamp 1636140361
transform 1 0 1363 0 1 5567
box 0 0 1 1
use contact_9  contact_9_43
timestamp 1636140361
transform 1 0 1359 0 1 5563
box 0 0 1 1
use contact_8  contact_8_49
timestamp 1636140361
transform 1 0 1360 0 1 5568
box 0 0 1 1
use contact_7  contact_7_50
timestamp 1636140361
transform 1 0 1363 0 1 5567
box 0 0 1 1
use contact_9  contact_9_50
timestamp 1636140361
transform 1 0 1359 0 1 5563
box 0 0 1 1
use contact_8  contact_8_56
timestamp 1636140361
transform 1 0 1360 0 1 5568
box 0 0 1 1
use pinv_20  pinv_20_21
timestamp 1636140361
transform 1 0 1472 0 -1 6720
box -36 -17 404 1177
use pinv_20  pinv_20_33
timestamp 1636140361
transform 1 0 0 0 1 6720
box -36 -17 404 1177
use pinv_20  pinv_20_32
timestamp 1636140361
transform 1 0 368 0 1 6720
box -36 -17 404 1177
use contact_9  contact_9_57
timestamp 1636140361
transform 1 0 163 0 1 6161
box 0 0 1 1
use contact_8  contact_8_59
timestamp 1636140361
transform 1 0 49 0 1 6166
box 0 0 1 1
use contact_7  contact_7_58
timestamp 1636140361
transform 1 0 167 0 1 6165
box 0 0 1 1
use contact_8  contact_8_58
timestamp 1636140361
transform 1 0 164 0 1 6166
box 0 0 1 1
use contact_7  contact_7_57
timestamp 1636140361
transform 1 0 52 0 1 6165
box 0 0 1 1
use contact_9  contact_9_51
timestamp 1636140361
transform 1 0 784 0 1 6161
box 0 0 1 1
use contact_8  contact_8_57
timestamp 1636140361
transform 1 0 785 0 1 6166
box 0 0 1 1
use contact_7  contact_7_65
timestamp 1636140361
transform 1 0 788 0 1 6165
box 0 0 1 1
use contact_9  contact_9_60
timestamp 1636140361
transform 1 0 416 0 1 6161
box 0 0 1 1
use contact_8  contact_8_68
timestamp 1636140361
transform 1 0 417 0 1 6166
box 0 0 1 1
use contact_7  contact_7_67
timestamp 1636140361
transform 1 0 420 0 1 6165
box 0 0 1 1
use contact_9  contact_9_53
timestamp 1636140361
transform 1 0 623 0 1 6683
box 0 0 1 1
use contact_8  contact_8_60
timestamp 1636140361
transform 1 0 624 0 1 6688
box 0 0 1 1
use contact_7  contact_7_59
timestamp 1636140361
transform 1 0 627 0 1 6687
box 0 0 1 1
use contact_9  contact_9_59
timestamp 1636140361
transform 1 0 623 0 1 6683
box 0 0 1 1
use contact_8  contact_8_67
timestamp 1636140361
transform 1 0 624 0 1 6688
box 0 0 1 1
use contact_7  contact_7_66
timestamp 1636140361
transform 1 0 627 0 1 6687
box 0 0 1 1
use pinv_20  pinv_20_38
timestamp 1636140361
transform 1 0 736 0 1 6720
box -36 -17 404 1177
use pinv_20  pinv_20_35
timestamp 1636140361
transform 1 0 1104 0 1 6720
box -36 -17 404 1177
use contact_7  contact_7_54
timestamp 1636140361
transform 1 0 1156 0 1 6165
box 0 0 1 1
use contact_8  contact_8_52
timestamp 1636140361
transform 1 0 1153 0 1 6166
box 0 0 1 1
use contact_9  contact_9_46
timestamp 1636140361
transform 1 0 1152 0 1 6161
box 0 0 1 1
use contact_9  contact_9_45
timestamp 1636140361
transform 1 0 1520 0 1 6161
box 0 0 1 1
use contact_8  contact_8_51
timestamp 1636140361
transform 1 0 1521 0 1 6166
box 0 0 1 1
use contact_7  contact_7_53
timestamp 1636140361
transform 1 0 1524 0 1 6165
box 0 0 1 1
use contact_9  contact_9_47
timestamp 1636140361
transform 1 0 1359 0 1 6683
box 0 0 1 1
use contact_8  contact_8_53
timestamp 1636140361
transform 1 0 1360 0 1 6688
box 0 0 1 1
use contact_7  contact_7_55
timestamp 1636140361
transform 1 0 1363 0 1 6687
box 0 0 1 1
use contact_9  contact_9_49
timestamp 1636140361
transform 1 0 1359 0 1 6683
box 0 0 1 1
use contact_8  contact_8_55
timestamp 1636140361
transform 1 0 1360 0 1 6688
box 0 0 1 1
use contact_7  contact_7_56
timestamp 1636140361
transform 1 0 1363 0 1 6687
box 0 0 1 1
use pinv_20  pinv_20_34
timestamp 1636140361
transform 1 0 1472 0 1 6720
box -36 -17 404 1177
use pinv_20  pinv_20_25
timestamp 1636140361
transform 1 0 0 0 -1 8960
box -36 -17 404 1177
use pinv_20  pinv_20_24
timestamp 1636140361
transform 1 0 368 0 -1 8960
box -36 -17 404 1177
use contact_7  contact_7_64
timestamp 1636140361
transform 1 0 52 0 1 7209
box 0 0 1 1
use contact_8  contact_8_66
timestamp 1636140361
transform 1 0 49 0 1 7210
box 0 0 1 1
use contact_7  contact_7_63
timestamp 1636140361
transform 1 0 167 0 1 7209
box 0 0 1 1
use contact_8  contact_8_64
timestamp 1636140361
transform 1 0 164 0 1 7210
box 0 0 1 1
use contact_9  contact_9_56
timestamp 1636140361
transform 1 0 163 0 1 7205
box 0 0 1 1
use contact_9  contact_9_52
timestamp 1636140361
transform 1 0 784 0 1 7205
box 0 0 1 1
use contact_8  contact_8_61
timestamp 1636140361
transform 1 0 785 0 1 7210
box 0 0 1 1
use contact_7  contact_7_60
timestamp 1636140361
transform 1 0 788 0 1 7209
box 0 0 1 1
use contact_9  contact_9_54
timestamp 1636140361
transform 1 0 416 0 1 7205
box 0 0 1 1
use contact_8  contact_8_63
timestamp 1636140361
transform 1 0 417 0 1 7210
box 0 0 1 1
use contact_7  contact_7_62
timestamp 1636140361
transform 1 0 420 0 1 7209
box 0 0 1 1
use contact_9  contact_9_66
timestamp 1636140361
transform 1 0 623 0 1 7803
box 0 0 1 1
use contact_8  contact_8_74
timestamp 1636140361
transform 1 0 624 0 1 7808
box 0 0 1 1
use contact_7  contact_7_75
timestamp 1636140361
transform 1 0 627 0 1 7807
box 0 0 1 1
use contact_9  contact_9_67
timestamp 1636140361
transform 1 0 623 0 1 7803
box 0 0 1 1
use contact_8  contact_8_75
timestamp 1636140361
transform 1 0 624 0 1 7808
box 0 0 1 1
use contact_7  contact_7_76
timestamp 1636140361
transform 1 0 627 0 1 7807
box 0 0 1 1
use pinv_20  pinv_20_37
timestamp 1636140361
transform 1 0 736 0 -1 8960
box -36 -17 404 1177
use pinv_20  pinv_20_29
timestamp 1636140361
transform 1 0 1104 0 -1 8960
box -36 -17 404 1177
use contact_7  contact_7_52
timestamp 1636140361
transform 1 0 1156 0 1 7209
box 0 0 1 1
use contact_8  contact_8_50
timestamp 1636140361
transform 1 0 1153 0 1 7210
box 0 0 1 1
use contact_9  contact_9_44
timestamp 1636140361
transform 1 0 1152 0 1 7205
box 0 0 1 1
use contact_7  contact_7_51
timestamp 1636140361
transform 1 0 1524 0 1 7209
box 0 0 1 1
use contact_9  contact_9_48
timestamp 1636140361
transform 1 0 1520 0 1 7205
box 0 0 1 1
use contact_8  contact_8_54
timestamp 1636140361
transform 1 0 1521 0 1 7210
box 0 0 1 1
use contact_9  contact_9_75
timestamp 1636140361
transform 1 0 1359 0 1 7803
box 0 0 1 1
use contact_8  contact_8_86
timestamp 1636140361
transform 1 0 1360 0 1 7808
box 0 0 1 1
use contact_7  contact_7_86
timestamp 1636140361
transform 1 0 1363 0 1 7807
box 0 0 1 1
use contact_9  contact_9_76
timestamp 1636140361
transform 1 0 1359 0 1 7803
box 0 0 1 1
use contact_8  contact_8_87
timestamp 1636140361
transform 1 0 1360 0 1 7808
box 0 0 1 1
use contact_7  contact_7_87
timestamp 1636140361
transform 1 0 1363 0 1 7807
box 0 0 1 1
use pinv_20  pinv_20_28
timestamp 1636140361
transform 1 0 1472 0 -1 8960
box -36 -17 404 1177
use contact_7  contact_7_69
timestamp 1636140361
transform 1 0 52 0 1 8405
box 0 0 1 1
use contact_9  contact_9_71
timestamp 1636140361
transform 1 0 163 0 1 8401
box 0 0 1 1
use contact_8  contact_8_80
timestamp 1636140361
transform 1 0 164 0 1 8406
box 0 0 1 1
use contact_7  contact_7_81
timestamp 1636140361
transform 1 0 167 0 1 8405
box 0 0 1 1
use contact_8  contact_8_81
timestamp 1636140361
transform 1 0 49 0 1 8406
box 0 0 1 1
use contact_9  contact_9_68
timestamp 1636140361
transform 1 0 163 0 1 9445
box 0 0 1 1
use contact_8  contact_8_76
timestamp 1636140361
transform 1 0 164 0 1 9450
box 0 0 1 1
use contact_7  contact_7_77
timestamp 1636140361
transform 1 0 167 0 1 9449
box 0 0 1 1
use contact_8  contact_8_77
timestamp 1636140361
transform 1 0 49 0 1 9450
box 0 0 1 1
use contact_7  contact_7_78
timestamp 1636140361
transform 1 0 52 0 1 9449
box 0 0 1 1
use pinv_20  pinv_20_26
timestamp 1636140361
transform 1 0 0 0 1 8960
box -36 -17 404 1177
use pinv_20  pinv_20_27
timestamp 1636140361
transform 1 0 368 0 1 8960
box -36 -17 404 1177
use contact_9  contact_9_61
timestamp 1636140361
transform 1 0 623 0 1 8923
box 0 0 1 1
use contact_9  contact_9_62
timestamp 1636140361
transform 1 0 784 0 1 8401
box 0 0 1 1
use contact_8  contact_8_70
timestamp 1636140361
transform 1 0 785 0 1 8406
box 0 0 1 1
use contact_7  contact_7_71
timestamp 1636140361
transform 1 0 788 0 1 8405
box 0 0 1 1
use contact_9  contact_9_64
timestamp 1636140361
transform 1 0 416 0 1 8401
box 0 0 1 1
use contact_8  contact_8_72
timestamp 1636140361
transform 1 0 417 0 1 8406
box 0 0 1 1
use contact_7  contact_7_73
timestamp 1636140361
transform 1 0 420 0 1 8405
box 0 0 1 1
use contact_9  contact_9_65
timestamp 1636140361
transform 1 0 623 0 1 8923
box 0 0 1 1
use contact_7  contact_7_74
timestamp 1636140361
transform 1 0 627 0 1 8927
box 0 0 1 1
use contact_8  contact_8_73
timestamp 1636140361
transform 1 0 624 0 1 8928
box 0 0 1 1
use contact_7  contact_7_70
timestamp 1636140361
transform 1 0 627 0 1 8927
box 0 0 1 1
use contact_8  contact_8_69
timestamp 1636140361
transform 1 0 624 0 1 8928
box 0 0 1 1
use contact_7  contact_7_80
timestamp 1636140361
transform 1 0 420 0 1 9449
box 0 0 1 1
use contact_8  contact_8_79
timestamp 1636140361
transform 1 0 417 0 1 9450
box 0 0 1 1
use contact_9  contact_9_70
timestamp 1636140361
transform 1 0 416 0 1 9445
box 0 0 1 1
use contact_7  contact_7_79
timestamp 1636140361
transform 1 0 788 0 1 9449
box 0 0 1 1
use contact_8  contact_8_78
timestamp 1636140361
transform 1 0 785 0 1 9450
box 0 0 1 1
use contact_9  contact_9_69
timestamp 1636140361
transform 1 0 784 0 1 9445
box 0 0 1 1
use pinv_20  pinv_20_36
timestamp 1636140361
transform 1 0 736 0 1 8960
box -36 -17 404 1177
use pinv_20  pinv_20_31
timestamp 1636140361
transform 1 0 1104 0 1 8960
box -36 -17 404 1177
use contact_7  contact_7_91
timestamp 1636140361
transform 1 0 1156 0 1 8405
box 0 0 1 1
use contact_8  contact_8_91
timestamp 1636140361
transform 1 0 1153 0 1 8406
box 0 0 1 1
use contact_9  contact_9_80
timestamp 1636140361
transform 1 0 1152 0 1 8401
box 0 0 1 1
use contact_7  contact_7_89
timestamp 1636140361
transform 1 0 1156 0 1 9449
box 0 0 1 1
use contact_8  contact_8_89
timestamp 1636140361
transform 1 0 1153 0 1 9450
box 0 0 1 1
use contact_9  contact_9_78
timestamp 1636140361
transform 1 0 1152 0 1 9445
box 0 0 1 1
use contact_9  contact_9_72
timestamp 1636140361
transform 1 0 1359 0 1 8923
box 0 0 1 1
use contact_9  contact_9_74
timestamp 1636140361
transform 1 0 1359 0 1 8923
box 0 0 1 1
use contact_9  contact_9_79
timestamp 1636140361
transform 1 0 1520 0 1 8401
box 0 0 1 1
use contact_8  contact_8_90
timestamp 1636140361
transform 1 0 1521 0 1 8406
box 0 0 1 1
use contact_7  contact_7_90
timestamp 1636140361
transform 1 0 1524 0 1 8405
box 0 0 1 1
use contact_8  contact_8_82
timestamp 1636140361
transform 1 0 1521 0 1 9450
box 0 0 1 1
use contact_7  contact_7_82
timestamp 1636140361
transform 1 0 1524 0 1 9449
box 0 0 1 1
use contact_8  contact_8_83
timestamp 1636140361
transform 1 0 1360 0 1 8928
box 0 0 1 1
use contact_7  contact_7_83
timestamp 1636140361
transform 1 0 1363 0 1 8927
box 0 0 1 1
use contact_8  contact_8_85
timestamp 1636140361
transform 1 0 1360 0 1 8928
box 0 0 1 1
use contact_7  contact_7_85
timestamp 1636140361
transform 1 0 1363 0 1 8927
box 0 0 1 1
use contact_9  contact_9_77
timestamp 1636140361
transform 1 0 1520 0 1 9445
box 0 0 1 1
use contact_8  contact_8_88
timestamp 1636140361
transform 1 0 1521 0 1 9450
box 0 0 1 1
use contact_7  contact_7_88
timestamp 1636140361
transform 1 0 1524 0 1 9449
box 0 0 1 1
use pinv_20  pinv_20_30
timestamp 1636140361
transform 1 0 1472 0 1 8960
box -36 -17 404 1177
use contact_7  contact_7_72
timestamp 1636140361
transform 1 0 627 0 1 10047
box 0 0 1 1
use contact_8  contact_8_71
timestamp 1636140361
transform 1 0 624 0 1 10048
box 0 0 1 1
use contact_9  contact_9_63
timestamp 1636140361
transform 1 0 623 0 1 10043
box 0 0 1 1
use contact_7  contact_7_84
timestamp 1636140361
transform 1 0 1363 0 1 10047
box 0 0 1 1
use contact_8  contact_8_84
timestamp 1636140361
transform 1 0 1360 0 1 10048
box 0 0 1 1
use contact_9  contact_9_73
timestamp 1636140361
transform 1 0 1359 0 1 10043
box 0 0 1 1
<< labels >>
rlabel metal2 s 78 261 78 261 4 in
port 1 nsew
rlabel metal2 s 1637 4741 1637 4741 4 out
port 2 nsew
rlabel metal3 s 656 2240 656 2240 4 gnd
port 4 nsew
rlabel metal3 s 1392 4480 1392 4480 4 gnd
port 4 nsew
rlabel metal3 s 656 4480 656 4480 4 gnd
port 4 nsew
rlabel metal3 s 1392 2240 1392 2240 4 gnd
port 4 nsew
rlabel metal3 s 656 6720 656 6720 4 gnd
port 4 nsew
rlabel metal3 s 656 8960 656 8960 4 gnd
port 4 nsew
rlabel metal3 s 1392 0 1392 0 4 gnd
port 4 nsew
rlabel metal3 s 1392 6720 1392 6720 4 gnd
port 4 nsew
rlabel metal3 s 1392 8960 1392 8960 4 gnd
port 4 nsew
rlabel metal3 s 656 0 656 0 4 gnd
port 4 nsew
rlabel metal3 s 656 10080 656 10080 4 vdd
port 3 nsew
rlabel metal3 s 656 7840 656 7840 4 vdd
port 3 nsew
rlabel metal3 s 656 3360 656 3360 4 vdd
port 3 nsew
rlabel metal3 s 656 3360 656 3360 4 vdd
port 3 nsew
rlabel metal3 s 1392 3360 1392 3360 4 vdd
port 3 nsew
rlabel metal3 s 1392 3360 1392 3360 4 vdd
port 3 nsew
rlabel metal3 s 1392 7840 1392 7840 4 vdd
port 3 nsew
rlabel metal3 s 656 1120 656 1120 4 vdd
port 3 nsew
rlabel metal3 s 1392 1120 1392 1120 4 vdd
port 3 nsew
rlabel metal3 s 1392 1120 1392 1120 4 vdd
port 3 nsew
rlabel metal3 s 656 1120 656 1120 4 vdd
port 3 nsew
rlabel metal3 s 656 5600 656 5600 4 vdd
port 3 nsew
rlabel metal3 s 1392 5600 1392 5600 4 vdd
port 3 nsew
rlabel metal3 s 1392 10080 1392 10080 4 vdd
port 3 nsew
<< properties >>
string FIXED_BBOX 1359 -37 1425 0
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_END 4882276
string GDS_START 4854004
<< end >>
