module ldpc(clk, rst, L1,
L2,
L3,
L4,
L5,
L6,
L7,
L8,
L9,
L10,
L11,
L12,
L13,
L14,
L15,
L16,
L17,
L18,
L19,
L20,
L21,
L22,
L23,
L24,
L25,
L26,
L27,
L28,
L29,
L30,
L31,
L32,
L33,
L34,
L35,
L36,
L37,
L38,
L39,
L40,
L41,
L42,
L43,
L44,
L45,
L46,
L47,
L48,
L49,
L50,
L51,
L52,
L53,
L54,
L55,
L56,
L57,
L58,
L59,
L60,
L61,
L62,
L63,
L64,
L65,
L66,
L67,
L68,
L69,
L70,
L71,
L72,
L73,
L74,
L75,
L76,
L77,
L78,
L79,
L80,
L81,
L82,
L83,
L84,
L85,
L86,
L87,
L88,
L89,
L90,
L91,
L92,
L93,
L94,
L95,
L96,
L97,
L98,
L99,
L100,
L101,
L102,
L103,
L104,
L105,
L106,
L107,
L108,
L109,
L110,
L111,
L112,
L113,
L114,
L115,
L116,
L117,
L118,
L119,
L120,
L121,
L122,
L123,
L124,
L125,
L126,
L127,
L128,
L129,
L130,
L131,
L132,
L133,
L134,
L135,
L136,
L137,
L138,
L139,
L140,
L141,
L142,
L143,
L144,
L145,
L146,
L147,
L148,
L149,
L150,
L151,
L152,
L153,
L154,
L155,
L156,
L157,
L158,
L159,
L160,
L161,
L162,
L163,
L164,
L165,
L166,
L167,
L168,
L169,
L170,
L171,
L172,
L173,
L174,
L175,
L176,
L177,
L178,
L179,
L180,
L181,
L182,
L183,
L184,
L185,
L186,
L187,
L188,
L189,
L190,
L191,
L192,
L193,
L194,
L195,
L196,
L197,
L198,
L199,
L200,
L201,
L202,
L203,
L204,
L205,
L206,
L207,
L208,
L209,
L210,
L211,
L212,
L213,
L214,
L215,
L216,
L217,
L218,
L219,
L220,
L221,
L222,
L223,
L224,
L225,
L226,
L227,
L228,
L229,
L230,
L231,
L232,
L233,
L234,
L235,
L236,
L237,
L238,
L239,
L240,
L241,
L242,
L243,
L244,
L245,
L246,
L247,
L248,
L249,
L250,
L251,
L252,
L253,
L254,
L255,
L256,
L257,
L258,
L259,
L260,
L261,
L262,
L263,
L264,
L265,
L266,
L267,
L268,
L269,
L270,
L271,
L272,
L273,
L274,
L275,
L276,
L277,
L278,
L279,
L280,
L281,
L282,
L283,
L284,
L285,
L286,
L287,
L288,
L289,
L290,
L291,
L292,
L293,
L294,
L295,
L296,
L297,
L298,
L299,
L300,
L301,
L302,
L303,
L304,
L305,
L306,
L307,
L308,
L309,
L310,
L311,
L312,
L313,
L314,
L315,
L316,
L317,
L318,
L319,
L320,
L321,
L322,
L323,
L324,
L325,
L326,
L327,
L328,
L329,
L330,
L331,
L332,
L333,
L334,
L335,
L336,
L337,
L338,
L339,
L340,
L341,
L342,
L343,
L344,
L345,
L346,
L347,
L348,
L349,
L350,
L351,
L352,
L353,
L354,
L355,
L356,
L357,
L358,
L359,
L360,
L361,
L362,
L363,
L364,
L365,
L366,
L367,
L368,
L369,
L370,
L371,
L372,
L373,
L374,
L375,
L376,
L377,
L378,
L379,
L380,
L381,
L382,
L383,
L384,
L385,
L386,
L387,
L388,
L389,
L390,
L391,
L392,
L393,
L394,
L395,
L396,
L397,
L398,
L399,
L400,
L401,
L402,
L403,
L404,
L405,
L406,
L407,
L408,
L409,
L410,
L411,
L412,
L413,
L414,
L415,
L416,
L417,
L418,
L419,
L420,
L421,
L422,
L423,
L424,
L425,
L426,
L427,
L428,
L429,
L430,
L431,
L432,
L433,
L434,
L435,
L436,
L437,
L438,
L439,
L440,
L441,
L442,
L443,
L444,
L445,
L446,
L447,
L448,
L449,
L450,
L451,
L452,
L453,
L454,
L455,
L456,
L457,
L458,
L459,
L460,
L461,
L462,
L463,
L464,
L465,
L466,
L467,
L468,
L469,
L470,
L471,
L472,
L473,
L474,
L475,
L476,
L477,
L478,
L479,
L480,
L481,
L482,
L483,
L484,
L485,
L486,
L487,
L488,
L489,
L490,
L491,
L492,
L493,
L494,
L495,
L496,
L497,
L498,
L499,
L500,
L501,
L502,
L503,
L504,
L505,
L506,
L507,
L508,
L509,
L510,
L511,
L512,
L513,
L514,
L515,
L516,
L517,
L518,
L519,
L520,
L521,
L522,
L523,
L524,
L525,
L526,
L527,
L528,
L529,
L530,
L531,
L532,
L533,
L534,
L535,
L536,
L537,
L538,
L539,
L540,
L541,
L542,
L543,
L544,
L545,
L546,
L547,
L548,
L549,
L550,
L551,
L552,
L553,
L554,
L555,
L556,
L557,
L558,
L559,
L560,
L561,
L562,
L563,
L564,
L565,
L566,
L567,
L568,
L569,
L570,
L571,
L572,
L573,
L574,
L575,
L576,
P1,
P2,
P3,
P4,
P5,
P6,
P7,
P8,
P9,
P10,
P11,
P12,
P13,
P14,
P15,
P16,
P17,
P18,
P19,
P20,
P21,
P22,
P23,
P24,
P25,
P26,
P27,
P28,
P29,
P30,
P31,
P32,
P33,
P34,
P35,
P36,
P37,
P38,
P39,
P40,
P41,
P42,
P43,
P44,
P45,
P46,
P47,
P48,
P49,
P50,
P51,
P52,
P53,
P54,
P55,
P56,
P57,
P58,
P59,
P60,
P61,
P62,
P63,
P64,
P65,
P66,
P67,
P68,
P69,
P70,
P71,
P72,
P73,
P74,
P75,
P76,
P77,
P78,
P79,
P80,
P81,
P82,
P83,
P84,
P85,
P86,
P87,
P88,
P89,
P90,
P91,
P92,
P93,
P94,
P95,
P96,
P97,
P98,
P99,
P100,
P101,
P102,
P103,
P104,
P105,
P106,
P107,
P108,
P109,
P110,
P111,
P112,
P113,
P114,
P115,
P116,
P117,
P118,
P119,
P120,
P121,
P122,
P123,
P124,
P125,
P126,
P127,
P128,
P129,
P130,
P131,
P132,
P133,
P134,
P135,
P136,
P137,
P138,
P139,
P140,
P141,
P142,
P143,
P144,
P145,
P146,
P147,
P148,
P149,
P150,
P151,
P152,
P153,
P154,
P155,
P156,
P157,
P158,
P159,
P160,
P161,
P162,
P163,
P164,
P165,
P166,
P167,
P168,
P169,
P170,
P171,
P172,
P173,
P174,
P175,
P176,
P177,
P178,
P179,
P180,
P181,
P182,
P183,
P184,
P185,
P186,
P187,
P188,
P189,
P190,
P191,
P192,
P193,
P194,
P195,
P196,
P197,
P198,
P199,
P200,
P201,
P202,
P203,
P204,
P205,
P206,
P207,
P208,
P209,
P210,
P211,
P212,
P213,
P214,
P215,
P216,
P217,
P218,
P219,
P220,
P221,
P222,
P223,
P224,
P225,
P226,
P227,
P228,
P229,
P230,
P231,
P232,
P233,
P234,
P235,
P236,
P237,
P238,
P239,
P240,
P241,
P242,
P243,
P244,
P245,
P246,
P247,
P248,
P249,
P250,
P251,
P252,
P253,
P254,
P255,
P256,
P257,
P258,
P259,
P260,
P261,
P262,
P263,
P264,
P265,
P266,
P267,
P268,
P269,
P270,
P271,
P272,
P273,
P274,
P275,
P276,
P277,
P278,
P279,
P280,
P281,
P282,
P283,
P284,
P285,
P286,
P287,
P288,
P289,
P290,
P291,
P292,
P293,
P294,
P295,
P296,
P297,
P298,
P299,
P300,
P301,
P302,
P303,
P304,
P305,
P306,
P307,
P308,
P309,
P310,
P311,
P312,
P313,
P314,
P315,
P316,
P317,
P318,
P319,
P320,
P321,
P322,
P323,
P324,
P325,
P326,
P327,
P328,
P329,
P330,
P331,
P332,
P333,
P334,
P335,
P336,
P337,
P338,
P339,
P340,
P341,
P342,
P343,
P344,
P345,
P346,
P347,
P348,
P349,
P350,
P351,
P352,
P353,
P354,
P355,
P356,
P357,
P358,
P359,
P360,
P361,
P362,
P363,
P364,
P365,
P366,
P367,
P368,
P369,
P370,
P371,
P372,
P373,
P374,
P375,
P376,
P377,
P378,
P379,
P380,
P381,
P382,
P383,
P384,
P385,
P386,
P387,
P388,
P389,
P390,
P391,
P392,
P393,
P394,
P395,
P396,
P397,
P398,
P399,
P400,
P401,
P402,
P403,
P404,
P405,
P406,
P407,
P408,
P409,
P410,
P411,
P412,
P413,
P414,
P415,
P416,
P417,
P418,
P419,
P420,
P421,
P422,
P423,
P424,
P425,
P426,
P427,
P428,
P429,
P430,
P431,
P432,
P433,
P434,
P435,
P436,
P437,
P438,
P439,
P440,
P441,
P442,
P443,
P444,
P445,
P446,
P447,
P448,
P449,
P450,
P451,
P452,
P453,
P454,
P455,
P456,
P457,
P458,
P459,
P460,
P461,
P462,
P463,
P464,
P465,
P466,
P467,
P468,
P469,
P470,
P471,
P472,
P473,
P474,
P475,
P476,
P477,
P478,
P479,
P480,
P481,
P482,
P483,
P484,
P485,
P486,
P487,
P488,
P489,
P490,
P491,
P492,
P493,
P494,
P495,
P496,
P497,
P498,
P499,
P500,
P501,
P502,
P503,
P504,
P505,
P506,
P507,
P508,
P509,
P510,
P511,
P512,
P513,
P514,
P515,
P516,
P517,
P518,
P519,
P520,
P521,
P522,
P523,
P524,
P525,
P526,
P527,
P528,
P529,
P530,
P531,
P532,
P533,
P534,
P535,
P536,
P537,
P538,
P539,
P540,
P541,
P542,
P543,
P544,
P545,
P546,
P547,
P548,
P549,
P550,
P551,
P552,
P553,
P554,
P555,
P556,
P557,
P558,
P559,
P560,
P561,
P562,
P563,
P564,
P565,
P566,
P567,
P568,
P569,
P570,
P571,
P572,
P573,
P574,
P575,
P576
);
input clk;
input rst;
input signed [31:0] L1;
input signed [31:0] L2;
input signed [31:0] L3;
input signed [31:0] L4;
input signed [31:0] L5;
input signed [31:0] L6;
input signed [31:0] L7;
input signed [31:0] L8;
input signed [31:0] L9;
input signed [31:0] L10;
input signed [31:0] L11;
input signed [31:0] L12;
input signed [31:0] L13;
input signed [31:0] L14;
input signed [31:0] L15;
input signed [31:0] L16;
input signed [31:0] L17;
input signed [31:0] L18;
input signed [31:0] L19;
input signed [31:0] L20;
input signed [31:0] L21;
input signed [31:0] L22;
input signed [31:0] L23;
input signed [31:0] L24;
input signed [31:0] L25;
input signed [31:0] L26;
input signed [31:0] L27;
input signed [31:0] L28;
input signed [31:0] L29;
input signed [31:0] L30;
input signed [31:0] L31;
input signed [31:0] L32;
input signed [31:0] L33;
input signed [31:0] L34;
input signed [31:0] L35;
input signed [31:0] L36;
input signed [31:0] L37;
input signed [31:0] L38;
input signed [31:0] L39;
input signed [31:0] L40;
input signed [31:0] L41;
input signed [31:0] L42;
input signed [31:0] L43;
input signed [31:0] L44;
input signed [31:0] L45;
input signed [31:0] L46;
input signed [31:0] L47;
input signed [31:0] L48;
input signed [31:0] L49;
input signed [31:0] L50;
input signed [31:0] L51;
input signed [31:0] L52;
input signed [31:0] L53;
input signed [31:0] L54;
input signed [31:0] L55;
input signed [31:0] L56;
input signed [31:0] L57;
input signed [31:0] L58;
input signed [31:0] L59;
input signed [31:0] L60;
input signed [31:0] L61;
input signed [31:0] L62;
input signed [31:0] L63;
input signed [31:0] L64;
input signed [31:0] L65;
input signed [31:0] L66;
input signed [31:0] L67;
input signed [31:0] L68;
input signed [31:0] L69;
input signed [31:0] L70;
input signed [31:0] L71;
input signed [31:0] L72;
input signed [31:0] L73;
input signed [31:0] L74;
input signed [31:0] L75;
input signed [31:0] L76;
input signed [31:0] L77;
input signed [31:0] L78;
input signed [31:0] L79;
input signed [31:0] L80;
input signed [31:0] L81;
input signed [31:0] L82;
input signed [31:0] L83;
input signed [31:0] L84;
input signed [31:0] L85;
input signed [31:0] L86;
input signed [31:0] L87;
input signed [31:0] L88;
input signed [31:0] L89;
input signed [31:0] L90;
input signed [31:0] L91;
input signed [31:0] L92;
input signed [31:0] L93;
input signed [31:0] L94;
input signed [31:0] L95;
input signed [31:0] L96;
input signed [31:0] L97;
input signed [31:0] L98;
input signed [31:0] L99;
input signed [31:0] L100;
input signed [31:0] L101;
input signed [31:0] L102;
input signed [31:0] L103;
input signed [31:0] L104;
input signed [31:0] L105;
input signed [31:0] L106;
input signed [31:0] L107;
input signed [31:0] L108;
input signed [31:0] L109;
input signed [31:0] L110;
input signed [31:0] L111;
input signed [31:0] L112;
input signed [31:0] L113;
input signed [31:0] L114;
input signed [31:0] L115;
input signed [31:0] L116;
input signed [31:0] L117;
input signed [31:0] L118;
input signed [31:0] L119;
input signed [31:0] L120;
input signed [31:0] L121;
input signed [31:0] L122;
input signed [31:0] L123;
input signed [31:0] L124;
input signed [31:0] L125;
input signed [31:0] L126;
input signed [31:0] L127;
input signed [31:0] L128;
input signed [31:0] L129;
input signed [31:0] L130;
input signed [31:0] L131;
input signed [31:0] L132;
input signed [31:0] L133;
input signed [31:0] L134;
input signed [31:0] L135;
input signed [31:0] L136;
input signed [31:0] L137;
input signed [31:0] L138;
input signed [31:0] L139;
input signed [31:0] L140;
input signed [31:0] L141;
input signed [31:0] L142;
input signed [31:0] L143;
input signed [31:0] L144;
input signed [31:0] L145;
input signed [31:0] L146;
input signed [31:0] L147;
input signed [31:0] L148;
input signed [31:0] L149;
input signed [31:0] L150;
input signed [31:0] L151;
input signed [31:0] L152;
input signed [31:0] L153;
input signed [31:0] L154;
input signed [31:0] L155;
input signed [31:0] L156;
input signed [31:0] L157;
input signed [31:0] L158;
input signed [31:0] L159;
input signed [31:0] L160;
input signed [31:0] L161;
input signed [31:0] L162;
input signed [31:0] L163;
input signed [31:0] L164;
input signed [31:0] L165;
input signed [31:0] L166;
input signed [31:0] L167;
input signed [31:0] L168;
input signed [31:0] L169;
input signed [31:0] L170;
input signed [31:0] L171;
input signed [31:0] L172;
input signed [31:0] L173;
input signed [31:0] L174;
input signed [31:0] L175;
input signed [31:0] L176;
input signed [31:0] L177;
input signed [31:0] L178;
input signed [31:0] L179;
input signed [31:0] L180;
input signed [31:0] L181;
input signed [31:0] L182;
input signed [31:0] L183;
input signed [31:0] L184;
input signed [31:0] L185;
input signed [31:0] L186;
input signed [31:0] L187;
input signed [31:0] L188;
input signed [31:0] L189;
input signed [31:0] L190;
input signed [31:0] L191;
input signed [31:0] L192;
input signed [31:0] L193;
input signed [31:0] L194;
input signed [31:0] L195;
input signed [31:0] L196;
input signed [31:0] L197;
input signed [31:0] L198;
input signed [31:0] L199;
input signed [31:0] L200;
input signed [31:0] L201;
input signed [31:0] L202;
input signed [31:0] L203;
input signed [31:0] L204;
input signed [31:0] L205;
input signed [31:0] L206;
input signed [31:0] L207;
input signed [31:0] L208;
input signed [31:0] L209;
input signed [31:0] L210;
input signed [31:0] L211;
input signed [31:0] L212;
input signed [31:0] L213;
input signed [31:0] L214;
input signed [31:0] L215;
input signed [31:0] L216;
input signed [31:0] L217;
input signed [31:0] L218;
input signed [31:0] L219;
input signed [31:0] L220;
input signed [31:0] L221;
input signed [31:0] L222;
input signed [31:0] L223;
input signed [31:0] L224;
input signed [31:0] L225;
input signed [31:0] L226;
input signed [31:0] L227;
input signed [31:0] L228;
input signed [31:0] L229;
input signed [31:0] L230;
input signed [31:0] L231;
input signed [31:0] L232;
input signed [31:0] L233;
input signed [31:0] L234;
input signed [31:0] L235;
input signed [31:0] L236;
input signed [31:0] L237;
input signed [31:0] L238;
input signed [31:0] L239;
input signed [31:0] L240;
input signed [31:0] L241;
input signed [31:0] L242;
input signed [31:0] L243;
input signed [31:0] L244;
input signed [31:0] L245;
input signed [31:0] L246;
input signed [31:0] L247;
input signed [31:0] L248;
input signed [31:0] L249;
input signed [31:0] L250;
input signed [31:0] L251;
input signed [31:0] L252;
input signed [31:0] L253;
input signed [31:0] L254;
input signed [31:0] L255;
input signed [31:0] L256;
input signed [31:0] L257;
input signed [31:0] L258;
input signed [31:0] L259;
input signed [31:0] L260;
input signed [31:0] L261;
input signed [31:0] L262;
input signed [31:0] L263;
input signed [31:0] L264;
input signed [31:0] L265;
input signed [31:0] L266;
input signed [31:0] L267;
input signed [31:0] L268;
input signed [31:0] L269;
input signed [31:0] L270;
input signed [31:0] L271;
input signed [31:0] L272;
input signed [31:0] L273;
input signed [31:0] L274;
input signed [31:0] L275;
input signed [31:0] L276;
input signed [31:0] L277;
input signed [31:0] L278;
input signed [31:0] L279;
input signed [31:0] L280;
input signed [31:0] L281;
input signed [31:0] L282;
input signed [31:0] L283;
input signed [31:0] L284;
input signed [31:0] L285;
input signed [31:0] L286;
input signed [31:0] L287;
input signed [31:0] L288;
input signed [31:0] L289;
input signed [31:0] L290;
input signed [31:0] L291;
input signed [31:0] L292;
input signed [31:0] L293;
input signed [31:0] L294;
input signed [31:0] L295;
input signed [31:0] L296;
input signed [31:0] L297;
input signed [31:0] L298;
input signed [31:0] L299;
input signed [31:0] L300;
input signed [31:0] L301;
input signed [31:0] L302;
input signed [31:0] L303;
input signed [31:0] L304;
input signed [31:0] L305;
input signed [31:0] L306;
input signed [31:0] L307;
input signed [31:0] L308;
input signed [31:0] L309;
input signed [31:0] L310;
input signed [31:0] L311;
input signed [31:0] L312;
input signed [31:0] L313;
input signed [31:0] L314;
input signed [31:0] L315;
input signed [31:0] L316;
input signed [31:0] L317;
input signed [31:0] L318;
input signed [31:0] L319;
input signed [31:0] L320;
input signed [31:0] L321;
input signed [31:0] L322;
input signed [31:0] L323;
input signed [31:0] L324;
input signed [31:0] L325;
input signed [31:0] L326;
input signed [31:0] L327;
input signed [31:0] L328;
input signed [31:0] L329;
input signed [31:0] L330;
input signed [31:0] L331;
input signed [31:0] L332;
input signed [31:0] L333;
input signed [31:0] L334;
input signed [31:0] L335;
input signed [31:0] L336;
input signed [31:0] L337;
input signed [31:0] L338;
input signed [31:0] L339;
input signed [31:0] L340;
input signed [31:0] L341;
input signed [31:0] L342;
input signed [31:0] L343;
input signed [31:0] L344;
input signed [31:0] L345;
input signed [31:0] L346;
input signed [31:0] L347;
input signed [31:0] L348;
input signed [31:0] L349;
input signed [31:0] L350;
input signed [31:0] L351;
input signed [31:0] L352;
input signed [31:0] L353;
input signed [31:0] L354;
input signed [31:0] L355;
input signed [31:0] L356;
input signed [31:0] L357;
input signed [31:0] L358;
input signed [31:0] L359;
input signed [31:0] L360;
input signed [31:0] L361;
input signed [31:0] L362;
input signed [31:0] L363;
input signed [31:0] L364;
input signed [31:0] L365;
input signed [31:0] L366;
input signed [31:0] L367;
input signed [31:0] L368;
input signed [31:0] L369;
input signed [31:0] L370;
input signed [31:0] L371;
input signed [31:0] L372;
input signed [31:0] L373;
input signed [31:0] L374;
input signed [31:0] L375;
input signed [31:0] L376;
input signed [31:0] L377;
input signed [31:0] L378;
input signed [31:0] L379;
input signed [31:0] L380;
input signed [31:0] L381;
input signed [31:0] L382;
input signed [31:0] L383;
input signed [31:0] L384;
input signed [31:0] L385;
input signed [31:0] L386;
input signed [31:0] L387;
input signed [31:0] L388;
input signed [31:0] L389;
input signed [31:0] L390;
input signed [31:0] L391;
input signed [31:0] L392;
input signed [31:0] L393;
input signed [31:0] L394;
input signed [31:0] L395;
input signed [31:0] L396;
input signed [31:0] L397;
input signed [31:0] L398;
input signed [31:0] L399;
input signed [31:0] L400;
input signed [31:0] L401;
input signed [31:0] L402;
input signed [31:0] L403;
input signed [31:0] L404;
input signed [31:0] L405;
input signed [31:0] L406;
input signed [31:0] L407;
input signed [31:0] L408;
input signed [31:0] L409;
input signed [31:0] L410;
input signed [31:0] L411;
input signed [31:0] L412;
input signed [31:0] L413;
input signed [31:0] L414;
input signed [31:0] L415;
input signed [31:0] L416;
input signed [31:0] L417;
input signed [31:0] L418;
input signed [31:0] L419;
input signed [31:0] L420;
input signed [31:0] L421;
input signed [31:0] L422;
input signed [31:0] L423;
input signed [31:0] L424;
input signed [31:0] L425;
input signed [31:0] L426;
input signed [31:0] L427;
input signed [31:0] L428;
input signed [31:0] L429;
input signed [31:0] L430;
input signed [31:0] L431;
input signed [31:0] L432;
input signed [31:0] L433;
input signed [31:0] L434;
input signed [31:0] L435;
input signed [31:0] L436;
input signed [31:0] L437;
input signed [31:0] L438;
input signed [31:0] L439;
input signed [31:0] L440;
input signed [31:0] L441;
input signed [31:0] L442;
input signed [31:0] L443;
input signed [31:0] L444;
input signed [31:0] L445;
input signed [31:0] L446;
input signed [31:0] L447;
input signed [31:0] L448;
input signed [31:0] L449;
input signed [31:0] L450;
input signed [31:0] L451;
input signed [31:0] L452;
input signed [31:0] L453;
input signed [31:0] L454;
input signed [31:0] L455;
input signed [31:0] L456;
input signed [31:0] L457;
input signed [31:0] L458;
input signed [31:0] L459;
input signed [31:0] L460;
input signed [31:0] L461;
input signed [31:0] L462;
input signed [31:0] L463;
input signed [31:0] L464;
input signed [31:0] L465;
input signed [31:0] L466;
input signed [31:0] L467;
input signed [31:0] L468;
input signed [31:0] L469;
input signed [31:0] L470;
input signed [31:0] L471;
input signed [31:0] L472;
input signed [31:0] L473;
input signed [31:0] L474;
input signed [31:0] L475;
input signed [31:0] L476;
input signed [31:0] L477;
input signed [31:0] L478;
input signed [31:0] L479;
input signed [31:0] L480;
input signed [31:0] L481;
input signed [31:0] L482;
input signed [31:0] L483;
input signed [31:0] L484;
input signed [31:0] L485;
input signed [31:0] L486;
input signed [31:0] L487;
input signed [31:0] L488;
input signed [31:0] L489;
input signed [31:0] L490;
input signed [31:0] L491;
input signed [31:0] L492;
input signed [31:0] L493;
input signed [31:0] L494;
input signed [31:0] L495;
input signed [31:0] L496;
input signed [31:0] L497;
input signed [31:0] L498;
input signed [31:0] L499;
input signed [31:0] L500;
input signed [31:0] L501;
input signed [31:0] L502;
input signed [31:0] L503;
input signed [31:0] L504;
input signed [31:0] L505;
input signed [31:0] L506;
input signed [31:0] L507;
input signed [31:0] L508;
input signed [31:0] L509;
input signed [31:0] L510;
input signed [31:0] L511;
input signed [31:0] L512;
input signed [31:0] L513;
input signed [31:0] L514;
input signed [31:0] L515;
input signed [31:0] L516;
input signed [31:0] L517;
input signed [31:0] L518;
input signed [31:0] L519;
input signed [31:0] L520;
input signed [31:0] L521;
input signed [31:0] L522;
input signed [31:0] L523;
input signed [31:0] L524;
input signed [31:0] L525;
input signed [31:0] L526;
input signed [31:0] L527;
input signed [31:0] L528;
input signed [31:0] L529;
input signed [31:0] L530;
input signed [31:0] L531;
input signed [31:0] L532;
input signed [31:0] L533;
input signed [31:0] L534;
input signed [31:0] L535;
input signed [31:0] L536;
input signed [31:0] L537;
input signed [31:0] L538;
input signed [31:0] L539;
input signed [31:0] L540;
input signed [31:0] L541;
input signed [31:0] L542;
input signed [31:0] L543;
input signed [31:0] L544;
input signed [31:0] L545;
input signed [31:0] L546;
input signed [31:0] L547;
input signed [31:0] L548;
input signed [31:0] L549;
input signed [31:0] L550;
input signed [31:0] L551;
input signed [31:0] L552;
input signed [31:0] L553;
input signed [31:0] L554;
input signed [31:0] L555;
input signed [31:0] L556;
input signed [31:0] L557;
input signed [31:0] L558;
input signed [31:0] L559;
input signed [31:0] L560;
input signed [31:0] L561;
input signed [31:0] L562;
input signed [31:0] L563;
input signed [31:0] L564;
input signed [31:0] L565;
input signed [31:0] L566;
input signed [31:0] L567;
input signed [31:0] L568;
input signed [31:0] L569;
input signed [31:0] L570;
input signed [31:0] L571;
input signed [31:0] L572;
input signed [31:0] L573;
input signed [31:0] L574;
input signed [31:0] L575;
input signed [31:0] L576;
output P1;
output P2;
output P3;
output P4;
output P5;
output P6;
output P7;
output P8;
output P9;
output P10;
output P11;
output P12;
output P13;
output P14;
output P15;
output P16;
output P17;
output P18;
output P19;
output P20;
output P21;
output P22;
output P23;
output P24;
output P25;
output P26;
output P27;
output P28;
output P29;
output P30;
output P31;
output P32;
output P33;
output P34;
output P35;
output P36;
output P37;
output P38;
output P39;
output P40;
output P41;
output P42;
output P43;
output P44;
output P45;
output P46;
output P47;
output P48;
output P49;
output P50;
output P51;
output P52;
output P53;
output P54;
output P55;
output P56;
output P57;
output P58;
output P59;
output P60;
output P61;
output P62;
output P63;
output P64;
output P65;
output P66;
output P67;
output P68;
output P69;
output P70;
output P71;
output P72;
output P73;
output P74;
output P75;
output P76;
output P77;
output P78;
output P79;
output P80;
output P81;
output P82;
output P83;
output P84;
output P85;
output P86;
output P87;
output P88;
output P89;
output P90;
output P91;
output P92;
output P93;
output P94;
output P95;
output P96;
output P97;
output P98;
output P99;
output P100;
output P101;
output P102;
output P103;
output P104;
output P105;
output P106;
output P107;
output P108;
output P109;
output P110;
output P111;
output P112;
output P113;
output P114;
output P115;
output P116;
output P117;
output P118;
output P119;
output P120;
output P121;
output P122;
output P123;
output P124;
output P125;
output P126;
output P127;
output P128;
output P129;
output P130;
output P131;
output P132;
output P133;
output P134;
output P135;
output P136;
output P137;
output P138;
output P139;
output P140;
output P141;
output P142;
output P143;
output P144;
output P145;
output P146;
output P147;
output P148;
output P149;
output P150;
output P151;
output P152;
output P153;
output P154;
output P155;
output P156;
output P157;
output P158;
output P159;
output P160;
output P161;
output P162;
output P163;
output P164;
output P165;
output P166;
output P167;
output P168;
output P169;
output P170;
output P171;
output P172;
output P173;
output P174;
output P175;
output P176;
output P177;
output P178;
output P179;
output P180;
output P181;
output P182;
output P183;
output P184;
output P185;
output P186;
output P187;
output P188;
output P189;
output P190;
output P191;
output P192;
output P193;
output P194;
output P195;
output P196;
output P197;
output P198;
output P199;
output P200;
output P201;
output P202;
output P203;
output P204;
output P205;
output P206;
output P207;
output P208;
output P209;
output P210;
output P211;
output P212;
output P213;
output P214;
output P215;
output P216;
output P217;
output P218;
output P219;
output P220;
output P221;
output P222;
output P223;
output P224;
output P225;
output P226;
output P227;
output P228;
output P229;
output P230;
output P231;
output P232;
output P233;
output P234;
output P235;
output P236;
output P237;
output P238;
output P239;
output P240;
output P241;
output P242;
output P243;
output P244;
output P245;
output P246;
output P247;
output P248;
output P249;
output P250;
output P251;
output P252;
output P253;
output P254;
output P255;
output P256;
output P257;
output P258;
output P259;
output P260;
output P261;
output P262;
output P263;
output P264;
output P265;
output P266;
output P267;
output P268;
output P269;
output P270;
output P271;
output P272;
output P273;
output P274;
output P275;
output P276;
output P277;
output P278;
output P279;
output P280;
output P281;
output P282;
output P283;
output P284;
output P285;
output P286;
output P287;
output P288;
output P289;
output P290;
output P291;
output P292;
output P293;
output P294;
output P295;
output P296;
output P297;
output P298;
output P299;
output P300;
output P301;
output P302;
output P303;
output P304;
output P305;
output P306;
output P307;
output P308;
output P309;
output P310;
output P311;
output P312;
output P313;
output P314;
output P315;
output P316;
output P317;
output P318;
output P319;
output P320;
output P321;
output P322;
output P323;
output P324;
output P325;
output P326;
output P327;
output P328;
output P329;
output P330;
output P331;
output P332;
output P333;
output P334;
output P335;
output P336;
output P337;
output P338;
output P339;
output P340;
output P341;
output P342;
output P343;
output P344;
output P345;
output P346;
output P347;
output P348;
output P349;
output P350;
output P351;
output P352;
output P353;
output P354;
output P355;
output P356;
output P357;
output P358;
output P359;
output P360;
output P361;
output P362;
output P363;
output P364;
output P365;
output P366;
output P367;
output P368;
output P369;
output P370;
output P371;
output P372;
output P373;
output P374;
output P375;
output P376;
output P377;
output P378;
output P379;
output P380;
output P381;
output P382;
output P383;
output P384;
output P385;
output P386;
output P387;
output P388;
output P389;
output P390;
output P391;
output P392;
output P393;
output P394;
output P395;
output P396;
output P397;
output P398;
output P399;
output P400;
output P401;
output P402;
output P403;
output P404;
output P405;
output P406;
output P407;
output P408;
output P409;
output P410;
output P411;
output P412;
output P413;
output P414;
output P415;
output P416;
output P417;
output P418;
output P419;
output P420;
output P421;
output P422;
output P423;
output P424;
output P425;
output P426;
output P427;
output P428;
output P429;
output P430;
output P431;
output P432;
output P433;
output P434;
output P435;
output P436;
output P437;
output P438;
output P439;
output P440;
output P441;
output P442;
output P443;
output P444;
output P445;
output P446;
output P447;
output P448;
output P449;
output P450;
output P451;
output P452;
output P453;
output P454;
output P455;
output P456;
output P457;
output P458;
output P459;
output P460;
output P461;
output P462;
output P463;
output P464;
output P465;
output P466;
output P467;
output P468;
output P469;
output P470;
output P471;
output P472;
output P473;
output P474;
output P475;
output P476;
output P477;
output P478;
output P479;
output P480;
output P481;
output P482;
output P483;
output P484;
output P485;
output P486;
output P487;
output P488;
output P489;
output P490;
output P491;
output P492;
output P493;
output P494;
output P495;
output P496;
output P497;
output P498;
output P499;
output P500;
output P501;
output P502;
output P503;
output P504;
output P505;
output P506;
output P507;
output P508;
output P509;
output P510;
output P511;
output P512;
output P513;
output P514;
output P515;
output P516;
output P517;
output P518;
output P519;
output P520;
output P521;
output P522;
output P523;
output P524;
output P525;
output P526;
output P527;
output P528;
output P529;
output P530;
output P531;
output P532;
output P533;
output P534;
output P535;
output P536;
output P537;
output P538;
output P539;
output P540;
output P541;
output P542;
output P543;
output P544;
output P545;
output P546;
output P547;
output P548;
output P549;
output P550;
output P551;
output P552;
output P553;
output P554;
output P555;
output P556;
output P557;
output P558;
output P559;
output P560;
output P561;
output P562;
output P563;
output P564;
output P565;
output P566;
output P567;
output P568;
output P569;
output P570;
output P571;
output P572;
output P573;
output P574;
output P575;
output P576;
wire signed [31:0] R1_48;
wire signed [31:0] R1_67;
wire signed [31:0] R1_206;
wire signed [31:0] R1_237;
wire signed [31:0] R1_290;
wire signed [31:0] R1_313;
wire signed [31:0] R2_25;
wire signed [31:0] R2_68;
wire signed [31:0] R2_207;
wire signed [31:0] R2_238;
wire signed [31:0] R2_291;
wire signed [31:0] R2_314;
wire signed [31:0] R3_26;
wire signed [31:0] R3_69;
wire signed [31:0] R3_208;
wire signed [31:0] R3_239;
wire signed [31:0] R3_292;
wire signed [31:0] R3_315;
wire signed [31:0] R4_27;
wire signed [31:0] R4_70;
wire signed [31:0] R4_209;
wire signed [31:0] R4_240;
wire signed [31:0] R4_293;
wire signed [31:0] R4_316;
wire signed [31:0] R5_28;
wire signed [31:0] R5_71;
wire signed [31:0] R5_210;
wire signed [31:0] R5_217;
wire signed [31:0] R5_294;
wire signed [31:0] R5_317;
wire signed [31:0] R6_29;
wire signed [31:0] R6_72;
wire signed [31:0] R6_211;
wire signed [31:0] R6_218;
wire signed [31:0] R6_295;
wire signed [31:0] R6_318;
wire signed [31:0] R7_30;
wire signed [31:0] R7_49;
wire signed [31:0] R7_212;
wire signed [31:0] R7_219;
wire signed [31:0] R7_296;
wire signed [31:0] R7_319;
wire signed [31:0] R8_31;
wire signed [31:0] R8_50;
wire signed [31:0] R8_213;
wire signed [31:0] R8_220;
wire signed [31:0] R8_297;
wire signed [31:0] R8_320;
wire signed [31:0] R9_32;
wire signed [31:0] R9_51;
wire signed [31:0] R9_214;
wire signed [31:0] R9_221;
wire signed [31:0] R9_298;
wire signed [31:0] R9_321;
wire signed [31:0] R10_33;
wire signed [31:0] R10_52;
wire signed [31:0] R10_215;
wire signed [31:0] R10_222;
wire signed [31:0] R10_299;
wire signed [31:0] R10_322;
wire signed [31:0] R11_34;
wire signed [31:0] R11_53;
wire signed [31:0] R11_216;
wire signed [31:0] R11_223;
wire signed [31:0] R11_300;
wire signed [31:0] R11_323;
wire signed [31:0] R12_35;
wire signed [31:0] R12_54;
wire signed [31:0] R12_193;
wire signed [31:0] R12_224;
wire signed [31:0] R12_301;
wire signed [31:0] R12_324;
wire signed [31:0] R13_36;
wire signed [31:0] R13_55;
wire signed [31:0] R13_194;
wire signed [31:0] R13_225;
wire signed [31:0] R13_302;
wire signed [31:0] R13_325;
wire signed [31:0] R14_37;
wire signed [31:0] R14_56;
wire signed [31:0] R14_195;
wire signed [31:0] R14_226;
wire signed [31:0] R14_303;
wire signed [31:0] R14_326;
wire signed [31:0] R15_38;
wire signed [31:0] R15_57;
wire signed [31:0] R15_196;
wire signed [31:0] R15_227;
wire signed [31:0] R15_304;
wire signed [31:0] R15_327;
wire signed [31:0] R16_39;
wire signed [31:0] R16_58;
wire signed [31:0] R16_197;
wire signed [31:0] R16_228;
wire signed [31:0] R16_305;
wire signed [31:0] R16_328;
wire signed [31:0] R17_40;
wire signed [31:0] R17_59;
wire signed [31:0] R17_198;
wire signed [31:0] R17_229;
wire signed [31:0] R17_306;
wire signed [31:0] R17_329;
wire signed [31:0] R18_41;
wire signed [31:0] R18_60;
wire signed [31:0] R18_199;
wire signed [31:0] R18_230;
wire signed [31:0] R18_307;
wire signed [31:0] R18_330;
wire signed [31:0] R19_42;
wire signed [31:0] R19_61;
wire signed [31:0] R19_200;
wire signed [31:0] R19_231;
wire signed [31:0] R19_308;
wire signed [31:0] R19_331;
wire signed [31:0] R20_43;
wire signed [31:0] R20_62;
wire signed [31:0] R20_201;
wire signed [31:0] R20_232;
wire signed [31:0] R20_309;
wire signed [31:0] R20_332;
wire signed [31:0] R21_44;
wire signed [31:0] R21_63;
wire signed [31:0] R21_202;
wire signed [31:0] R21_233;
wire signed [31:0] R21_310;
wire signed [31:0] R21_333;
wire signed [31:0] R22_45;
wire signed [31:0] R22_64;
wire signed [31:0] R22_203;
wire signed [31:0] R22_234;
wire signed [31:0] R22_311;
wire signed [31:0] R22_334;
wire signed [31:0] R23_46;
wire signed [31:0] R23_65;
wire signed [31:0] R23_204;
wire signed [31:0] R23_235;
wire signed [31:0] R23_312;
wire signed [31:0] R23_335;
wire signed [31:0] R24_47;
wire signed [31:0] R24_66;
wire signed [31:0] R24_205;
wire signed [31:0] R24_236;
wire signed [31:0] R24_289;
wire signed [31:0] R24_336;
wire signed [31:0] R25_31;
wire signed [31:0] R25_126;
wire signed [31:0] R25_164;
wire signed [31:0] R25_171;
wire signed [31:0] R25_268;
wire signed [31:0] R25_313;
wire signed [31:0] R25_337;
wire signed [31:0] R26_32;
wire signed [31:0] R26_127;
wire signed [31:0] R26_165;
wire signed [31:0] R26_172;
wire signed [31:0] R26_269;
wire signed [31:0] R26_314;
wire signed [31:0] R26_338;
wire signed [31:0] R27_33;
wire signed [31:0] R27_128;
wire signed [31:0] R27_166;
wire signed [31:0] R27_173;
wire signed [31:0] R27_270;
wire signed [31:0] R27_315;
wire signed [31:0] R27_339;
wire signed [31:0] R28_34;
wire signed [31:0] R28_129;
wire signed [31:0] R28_167;
wire signed [31:0] R28_174;
wire signed [31:0] R28_271;
wire signed [31:0] R28_316;
wire signed [31:0] R28_340;
wire signed [31:0] R29_35;
wire signed [31:0] R29_130;
wire signed [31:0] R29_168;
wire signed [31:0] R29_175;
wire signed [31:0] R29_272;
wire signed [31:0] R29_317;
wire signed [31:0] R29_341;
wire signed [31:0] R30_36;
wire signed [31:0] R30_131;
wire signed [31:0] R30_145;
wire signed [31:0] R30_176;
wire signed [31:0] R30_273;
wire signed [31:0] R30_318;
wire signed [31:0] R30_342;
wire signed [31:0] R31_37;
wire signed [31:0] R31_132;
wire signed [31:0] R31_146;
wire signed [31:0] R31_177;
wire signed [31:0] R31_274;
wire signed [31:0] R31_319;
wire signed [31:0] R31_343;
wire signed [31:0] R32_38;
wire signed [31:0] R32_133;
wire signed [31:0] R32_147;
wire signed [31:0] R32_178;
wire signed [31:0] R32_275;
wire signed [31:0] R32_320;
wire signed [31:0] R32_344;
wire signed [31:0] R33_39;
wire signed [31:0] R33_134;
wire signed [31:0] R33_148;
wire signed [31:0] R33_179;
wire signed [31:0] R33_276;
wire signed [31:0] R33_321;
wire signed [31:0] R33_345;
wire signed [31:0] R34_40;
wire signed [31:0] R34_135;
wire signed [31:0] R34_149;
wire signed [31:0] R34_180;
wire signed [31:0] R34_277;
wire signed [31:0] R34_322;
wire signed [31:0] R34_346;
wire signed [31:0] R35_41;
wire signed [31:0] R35_136;
wire signed [31:0] R35_150;
wire signed [31:0] R35_181;
wire signed [31:0] R35_278;
wire signed [31:0] R35_323;
wire signed [31:0] R35_347;
wire signed [31:0] R36_42;
wire signed [31:0] R36_137;
wire signed [31:0] R36_151;
wire signed [31:0] R36_182;
wire signed [31:0] R36_279;
wire signed [31:0] R36_324;
wire signed [31:0] R36_348;
wire signed [31:0] R37_43;
wire signed [31:0] R37_138;
wire signed [31:0] R37_152;
wire signed [31:0] R37_183;
wire signed [31:0] R37_280;
wire signed [31:0] R37_325;
wire signed [31:0] R37_349;
wire signed [31:0] R38_44;
wire signed [31:0] R38_139;
wire signed [31:0] R38_153;
wire signed [31:0] R38_184;
wire signed [31:0] R38_281;
wire signed [31:0] R38_326;
wire signed [31:0] R38_350;
wire signed [31:0] R39_45;
wire signed [31:0] R39_140;
wire signed [31:0] R39_154;
wire signed [31:0] R39_185;
wire signed [31:0] R39_282;
wire signed [31:0] R39_327;
wire signed [31:0] R39_351;
wire signed [31:0] R40_46;
wire signed [31:0] R40_141;
wire signed [31:0] R40_155;
wire signed [31:0] R40_186;
wire signed [31:0] R40_283;
wire signed [31:0] R40_328;
wire signed [31:0] R40_352;
wire signed [31:0] R41_47;
wire signed [31:0] R41_142;
wire signed [31:0] R41_156;
wire signed [31:0] R41_187;
wire signed [31:0] R41_284;
wire signed [31:0] R41_329;
wire signed [31:0] R41_353;
wire signed [31:0] R42_48;
wire signed [31:0] R42_143;
wire signed [31:0] R42_157;
wire signed [31:0] R42_188;
wire signed [31:0] R42_285;
wire signed [31:0] R42_330;
wire signed [31:0] R42_354;
wire signed [31:0] R43_25;
wire signed [31:0] R43_144;
wire signed [31:0] R43_158;
wire signed [31:0] R43_189;
wire signed [31:0] R43_286;
wire signed [31:0] R43_331;
wire signed [31:0] R43_355;
wire signed [31:0] R44_26;
wire signed [31:0] R44_121;
wire signed [31:0] R44_159;
wire signed [31:0] R44_190;
wire signed [31:0] R44_287;
wire signed [31:0] R44_332;
wire signed [31:0] R44_356;
wire signed [31:0] R45_27;
wire signed [31:0] R45_122;
wire signed [31:0] R45_160;
wire signed [31:0] R45_191;
wire signed [31:0] R45_288;
wire signed [31:0] R45_333;
wire signed [31:0] R45_357;
wire signed [31:0] R46_28;
wire signed [31:0] R46_123;
wire signed [31:0] R46_161;
wire signed [31:0] R46_192;
wire signed [31:0] R46_265;
wire signed [31:0] R46_334;
wire signed [31:0] R46_358;
wire signed [31:0] R47_29;
wire signed [31:0] R47_124;
wire signed [31:0] R47_162;
wire signed [31:0] R47_169;
wire signed [31:0] R47_266;
wire signed [31:0] R47_335;
wire signed [31:0] R47_359;
wire signed [31:0] R48_30;
wire signed [31:0] R48_125;
wire signed [31:0] R48_163;
wire signed [31:0] R48_170;
wire signed [31:0] R48_267;
wire signed [31:0] R48_336;
wire signed [31:0] R48_360;
wire signed [31:0] R49_79;
wire signed [31:0] R49_102;
wire signed [31:0] R49_141;
wire signed [31:0] R49_177;
wire signed [31:0] R49_265;
wire signed [31:0] R49_337;
wire signed [31:0] R49_361;
wire signed [31:0] R50_80;
wire signed [31:0] R50_103;
wire signed [31:0] R50_142;
wire signed [31:0] R50_178;
wire signed [31:0] R50_266;
wire signed [31:0] R50_338;
wire signed [31:0] R50_362;
wire signed [31:0] R51_81;
wire signed [31:0] R51_104;
wire signed [31:0] R51_143;
wire signed [31:0] R51_179;
wire signed [31:0] R51_267;
wire signed [31:0] R51_339;
wire signed [31:0] R51_363;
wire signed [31:0] R52_82;
wire signed [31:0] R52_105;
wire signed [31:0] R52_144;
wire signed [31:0] R52_180;
wire signed [31:0] R52_268;
wire signed [31:0] R52_340;
wire signed [31:0] R52_364;
wire signed [31:0] R53_83;
wire signed [31:0] R53_106;
wire signed [31:0] R53_121;
wire signed [31:0] R53_181;
wire signed [31:0] R53_269;
wire signed [31:0] R53_341;
wire signed [31:0] R53_365;
wire signed [31:0] R54_84;
wire signed [31:0] R54_107;
wire signed [31:0] R54_122;
wire signed [31:0] R54_182;
wire signed [31:0] R54_270;
wire signed [31:0] R54_342;
wire signed [31:0] R54_366;
wire signed [31:0] R55_85;
wire signed [31:0] R55_108;
wire signed [31:0] R55_123;
wire signed [31:0] R55_183;
wire signed [31:0] R55_271;
wire signed [31:0] R55_343;
wire signed [31:0] R55_367;
wire signed [31:0] R56_86;
wire signed [31:0] R56_109;
wire signed [31:0] R56_124;
wire signed [31:0] R56_184;
wire signed [31:0] R56_272;
wire signed [31:0] R56_344;
wire signed [31:0] R56_368;
wire signed [31:0] R57_87;
wire signed [31:0] R57_110;
wire signed [31:0] R57_125;
wire signed [31:0] R57_185;
wire signed [31:0] R57_273;
wire signed [31:0] R57_345;
wire signed [31:0] R57_369;
wire signed [31:0] R58_88;
wire signed [31:0] R58_111;
wire signed [31:0] R58_126;
wire signed [31:0] R58_186;
wire signed [31:0] R58_274;
wire signed [31:0] R58_346;
wire signed [31:0] R58_370;
wire signed [31:0] R59_89;
wire signed [31:0] R59_112;
wire signed [31:0] R59_127;
wire signed [31:0] R59_187;
wire signed [31:0] R59_275;
wire signed [31:0] R59_347;
wire signed [31:0] R59_371;
wire signed [31:0] R60_90;
wire signed [31:0] R60_113;
wire signed [31:0] R60_128;
wire signed [31:0] R60_188;
wire signed [31:0] R60_276;
wire signed [31:0] R60_348;
wire signed [31:0] R60_372;
wire signed [31:0] R61_91;
wire signed [31:0] R61_114;
wire signed [31:0] R61_129;
wire signed [31:0] R61_189;
wire signed [31:0] R61_277;
wire signed [31:0] R61_349;
wire signed [31:0] R61_373;
wire signed [31:0] R62_92;
wire signed [31:0] R62_115;
wire signed [31:0] R62_130;
wire signed [31:0] R62_190;
wire signed [31:0] R62_278;
wire signed [31:0] R62_350;
wire signed [31:0] R62_374;
wire signed [31:0] R63_93;
wire signed [31:0] R63_116;
wire signed [31:0] R63_131;
wire signed [31:0] R63_191;
wire signed [31:0] R63_279;
wire signed [31:0] R63_351;
wire signed [31:0] R63_375;
wire signed [31:0] R64_94;
wire signed [31:0] R64_117;
wire signed [31:0] R64_132;
wire signed [31:0] R64_192;
wire signed [31:0] R64_280;
wire signed [31:0] R64_352;
wire signed [31:0] R64_376;
wire signed [31:0] R65_95;
wire signed [31:0] R65_118;
wire signed [31:0] R65_133;
wire signed [31:0] R65_169;
wire signed [31:0] R65_281;
wire signed [31:0] R65_353;
wire signed [31:0] R65_377;
wire signed [31:0] R66_96;
wire signed [31:0] R66_119;
wire signed [31:0] R66_134;
wire signed [31:0] R66_170;
wire signed [31:0] R66_282;
wire signed [31:0] R66_354;
wire signed [31:0] R66_378;
wire signed [31:0] R67_73;
wire signed [31:0] R67_120;
wire signed [31:0] R67_135;
wire signed [31:0] R67_171;
wire signed [31:0] R67_283;
wire signed [31:0] R67_355;
wire signed [31:0] R67_379;
wire signed [31:0] R68_74;
wire signed [31:0] R68_97;
wire signed [31:0] R68_136;
wire signed [31:0] R68_172;
wire signed [31:0] R68_284;
wire signed [31:0] R68_356;
wire signed [31:0] R68_380;
wire signed [31:0] R69_75;
wire signed [31:0] R69_98;
wire signed [31:0] R69_137;
wire signed [31:0] R69_173;
wire signed [31:0] R69_285;
wire signed [31:0] R69_357;
wire signed [31:0] R69_381;
wire signed [31:0] R70_76;
wire signed [31:0] R70_99;
wire signed [31:0] R70_138;
wire signed [31:0] R70_174;
wire signed [31:0] R70_286;
wire signed [31:0] R70_358;
wire signed [31:0] R70_382;
wire signed [31:0] R71_77;
wire signed [31:0] R71_100;
wire signed [31:0] R71_139;
wire signed [31:0] R71_175;
wire signed [31:0] R71_287;
wire signed [31:0] R71_359;
wire signed [31:0] R71_383;
wire signed [31:0] R72_78;
wire signed [31:0] R72_101;
wire signed [31:0] R72_140;
wire signed [31:0] R72_176;
wire signed [31:0] R72_288;
wire signed [31:0] R72_360;
wire signed [31:0] R72_384;
wire signed [31:0] R73_16;
wire signed [31:0] R73_60;
wire signed [31:0] R73_209;
wire signed [31:0] R73_223;
wire signed [31:0] R73_361;
wire signed [31:0] R73_385;
wire signed [31:0] R74_17;
wire signed [31:0] R74_61;
wire signed [31:0] R74_210;
wire signed [31:0] R74_224;
wire signed [31:0] R74_362;
wire signed [31:0] R74_386;
wire signed [31:0] R75_18;
wire signed [31:0] R75_62;
wire signed [31:0] R75_211;
wire signed [31:0] R75_225;
wire signed [31:0] R75_363;
wire signed [31:0] R75_387;
wire signed [31:0] R76_19;
wire signed [31:0] R76_63;
wire signed [31:0] R76_212;
wire signed [31:0] R76_226;
wire signed [31:0] R76_364;
wire signed [31:0] R76_388;
wire signed [31:0] R77_20;
wire signed [31:0] R77_64;
wire signed [31:0] R77_213;
wire signed [31:0] R77_227;
wire signed [31:0] R77_365;
wire signed [31:0] R77_389;
wire signed [31:0] R78_21;
wire signed [31:0] R78_65;
wire signed [31:0] R78_214;
wire signed [31:0] R78_228;
wire signed [31:0] R78_366;
wire signed [31:0] R78_390;
wire signed [31:0] R79_22;
wire signed [31:0] R79_66;
wire signed [31:0] R79_215;
wire signed [31:0] R79_229;
wire signed [31:0] R79_367;
wire signed [31:0] R79_391;
wire signed [31:0] R80_23;
wire signed [31:0] R80_67;
wire signed [31:0] R80_216;
wire signed [31:0] R80_230;
wire signed [31:0] R80_368;
wire signed [31:0] R80_392;
wire signed [31:0] R81_24;
wire signed [31:0] R81_68;
wire signed [31:0] R81_193;
wire signed [31:0] R81_231;
wire signed [31:0] R81_369;
wire signed [31:0] R81_393;
wire signed [31:0] R82_1;
wire signed [31:0] R82_69;
wire signed [31:0] R82_194;
wire signed [31:0] R82_232;
wire signed [31:0] R82_370;
wire signed [31:0] R82_394;
wire signed [31:0] R83_2;
wire signed [31:0] R83_70;
wire signed [31:0] R83_195;
wire signed [31:0] R83_233;
wire signed [31:0] R83_371;
wire signed [31:0] R83_395;
wire signed [31:0] R84_3;
wire signed [31:0] R84_71;
wire signed [31:0] R84_196;
wire signed [31:0] R84_234;
wire signed [31:0] R84_372;
wire signed [31:0] R84_396;
wire signed [31:0] R85_4;
wire signed [31:0] R85_72;
wire signed [31:0] R85_197;
wire signed [31:0] R85_235;
wire signed [31:0] R85_373;
wire signed [31:0] R85_397;
wire signed [31:0] R86_5;
wire signed [31:0] R86_49;
wire signed [31:0] R86_198;
wire signed [31:0] R86_236;
wire signed [31:0] R86_374;
wire signed [31:0] R86_398;
wire signed [31:0] R87_6;
wire signed [31:0] R87_50;
wire signed [31:0] R87_199;
wire signed [31:0] R87_237;
wire signed [31:0] R87_375;
wire signed [31:0] R87_399;
wire signed [31:0] R88_7;
wire signed [31:0] R88_51;
wire signed [31:0] R88_200;
wire signed [31:0] R88_238;
wire signed [31:0] R88_376;
wire signed [31:0] R88_400;
wire signed [31:0] R89_8;
wire signed [31:0] R89_52;
wire signed [31:0] R89_201;
wire signed [31:0] R89_239;
wire signed [31:0] R89_377;
wire signed [31:0] R89_401;
wire signed [31:0] R90_9;
wire signed [31:0] R90_53;
wire signed [31:0] R90_202;
wire signed [31:0] R90_240;
wire signed [31:0] R90_378;
wire signed [31:0] R90_402;
wire signed [31:0] R91_10;
wire signed [31:0] R91_54;
wire signed [31:0] R91_203;
wire signed [31:0] R91_217;
wire signed [31:0] R91_379;
wire signed [31:0] R91_403;
wire signed [31:0] R92_11;
wire signed [31:0] R92_55;
wire signed [31:0] R92_204;
wire signed [31:0] R92_218;
wire signed [31:0] R92_380;
wire signed [31:0] R92_404;
wire signed [31:0] R93_12;
wire signed [31:0] R93_56;
wire signed [31:0] R93_205;
wire signed [31:0] R93_219;
wire signed [31:0] R93_381;
wire signed [31:0] R93_405;
wire signed [31:0] R94_13;
wire signed [31:0] R94_57;
wire signed [31:0] R94_206;
wire signed [31:0] R94_220;
wire signed [31:0] R94_382;
wire signed [31:0] R94_406;
wire signed [31:0] R95_14;
wire signed [31:0] R95_58;
wire signed [31:0] R95_207;
wire signed [31:0] R95_221;
wire signed [31:0] R95_383;
wire signed [31:0] R95_407;
wire signed [31:0] R96_15;
wire signed [31:0] R96_59;
wire signed [31:0] R96_208;
wire signed [31:0] R96_222;
wire signed [31:0] R96_384;
wire signed [31:0] R96_408;
wire signed [31:0] R97_58;
wire signed [31:0] R97_166;
wire signed [31:0] R97_227;
wire signed [31:0] R97_259;
wire signed [31:0] R97_385;
wire signed [31:0] R97_409;
wire signed [31:0] R98_59;
wire signed [31:0] R98_167;
wire signed [31:0] R98_228;
wire signed [31:0] R98_260;
wire signed [31:0] R98_386;
wire signed [31:0] R98_410;
wire signed [31:0] R99_60;
wire signed [31:0] R99_168;
wire signed [31:0] R99_229;
wire signed [31:0] R99_261;
wire signed [31:0] R99_387;
wire signed [31:0] R99_411;
wire signed [31:0] R100_61;
wire signed [31:0] R100_145;
wire signed [31:0] R100_230;
wire signed [31:0] R100_262;
wire signed [31:0] R100_388;
wire signed [31:0] R100_412;
wire signed [31:0] R101_62;
wire signed [31:0] R101_146;
wire signed [31:0] R101_231;
wire signed [31:0] R101_263;
wire signed [31:0] R101_389;
wire signed [31:0] R101_413;
wire signed [31:0] R102_63;
wire signed [31:0] R102_147;
wire signed [31:0] R102_232;
wire signed [31:0] R102_264;
wire signed [31:0] R102_390;
wire signed [31:0] R102_414;
wire signed [31:0] R103_64;
wire signed [31:0] R103_148;
wire signed [31:0] R103_233;
wire signed [31:0] R103_241;
wire signed [31:0] R103_391;
wire signed [31:0] R103_415;
wire signed [31:0] R104_65;
wire signed [31:0] R104_149;
wire signed [31:0] R104_234;
wire signed [31:0] R104_242;
wire signed [31:0] R104_392;
wire signed [31:0] R104_416;
wire signed [31:0] R105_66;
wire signed [31:0] R105_150;
wire signed [31:0] R105_235;
wire signed [31:0] R105_243;
wire signed [31:0] R105_393;
wire signed [31:0] R105_417;
wire signed [31:0] R106_67;
wire signed [31:0] R106_151;
wire signed [31:0] R106_236;
wire signed [31:0] R106_244;
wire signed [31:0] R106_394;
wire signed [31:0] R106_418;
wire signed [31:0] R107_68;
wire signed [31:0] R107_152;
wire signed [31:0] R107_237;
wire signed [31:0] R107_245;
wire signed [31:0] R107_395;
wire signed [31:0] R107_419;
wire signed [31:0] R108_69;
wire signed [31:0] R108_153;
wire signed [31:0] R108_238;
wire signed [31:0] R108_246;
wire signed [31:0] R108_396;
wire signed [31:0] R108_420;
wire signed [31:0] R109_70;
wire signed [31:0] R109_154;
wire signed [31:0] R109_239;
wire signed [31:0] R109_247;
wire signed [31:0] R109_397;
wire signed [31:0] R109_421;
wire signed [31:0] R110_71;
wire signed [31:0] R110_155;
wire signed [31:0] R110_240;
wire signed [31:0] R110_248;
wire signed [31:0] R110_398;
wire signed [31:0] R110_422;
wire signed [31:0] R111_72;
wire signed [31:0] R111_156;
wire signed [31:0] R111_217;
wire signed [31:0] R111_249;
wire signed [31:0] R111_399;
wire signed [31:0] R111_423;
wire signed [31:0] R112_49;
wire signed [31:0] R112_157;
wire signed [31:0] R112_218;
wire signed [31:0] R112_250;
wire signed [31:0] R112_400;
wire signed [31:0] R112_424;
wire signed [31:0] R113_50;
wire signed [31:0] R113_158;
wire signed [31:0] R113_219;
wire signed [31:0] R113_251;
wire signed [31:0] R113_401;
wire signed [31:0] R113_425;
wire signed [31:0] R114_51;
wire signed [31:0] R114_159;
wire signed [31:0] R114_220;
wire signed [31:0] R114_252;
wire signed [31:0] R114_402;
wire signed [31:0] R114_426;
wire signed [31:0] R115_52;
wire signed [31:0] R115_160;
wire signed [31:0] R115_221;
wire signed [31:0] R115_253;
wire signed [31:0] R115_403;
wire signed [31:0] R115_427;
wire signed [31:0] R116_53;
wire signed [31:0] R116_161;
wire signed [31:0] R116_222;
wire signed [31:0] R116_254;
wire signed [31:0] R116_404;
wire signed [31:0] R116_428;
wire signed [31:0] R117_54;
wire signed [31:0] R117_162;
wire signed [31:0] R117_223;
wire signed [31:0] R117_255;
wire signed [31:0] R117_405;
wire signed [31:0] R117_429;
wire signed [31:0] R118_55;
wire signed [31:0] R118_163;
wire signed [31:0] R118_224;
wire signed [31:0] R118_256;
wire signed [31:0] R118_406;
wire signed [31:0] R118_430;
wire signed [31:0] R119_56;
wire signed [31:0] R119_164;
wire signed [31:0] R119_225;
wire signed [31:0] R119_257;
wire signed [31:0] R119_407;
wire signed [31:0] R119_431;
wire signed [31:0] R120_57;
wire signed [31:0] R120_165;
wire signed [31:0] R120_226;
wire signed [31:0] R120_258;
wire signed [31:0] R120_408;
wire signed [31:0] R120_432;
wire signed [31:0] R121_108;
wire signed [31:0] R121_131;
wire signed [31:0] R121_189;
wire signed [31:0] R121_284;
wire signed [31:0] R121_289;
wire signed [31:0] R121_409;
wire signed [31:0] R121_433;
wire signed [31:0] R122_109;
wire signed [31:0] R122_132;
wire signed [31:0] R122_190;
wire signed [31:0] R122_285;
wire signed [31:0] R122_290;
wire signed [31:0] R122_410;
wire signed [31:0] R122_434;
wire signed [31:0] R123_110;
wire signed [31:0] R123_133;
wire signed [31:0] R123_191;
wire signed [31:0] R123_286;
wire signed [31:0] R123_291;
wire signed [31:0] R123_411;
wire signed [31:0] R123_435;
wire signed [31:0] R124_111;
wire signed [31:0] R124_134;
wire signed [31:0] R124_192;
wire signed [31:0] R124_287;
wire signed [31:0] R124_292;
wire signed [31:0] R124_412;
wire signed [31:0] R124_436;
wire signed [31:0] R125_112;
wire signed [31:0] R125_135;
wire signed [31:0] R125_169;
wire signed [31:0] R125_288;
wire signed [31:0] R125_293;
wire signed [31:0] R125_413;
wire signed [31:0] R125_437;
wire signed [31:0] R126_113;
wire signed [31:0] R126_136;
wire signed [31:0] R126_170;
wire signed [31:0] R126_265;
wire signed [31:0] R126_294;
wire signed [31:0] R126_414;
wire signed [31:0] R126_438;
wire signed [31:0] R127_114;
wire signed [31:0] R127_137;
wire signed [31:0] R127_171;
wire signed [31:0] R127_266;
wire signed [31:0] R127_295;
wire signed [31:0] R127_415;
wire signed [31:0] R127_439;
wire signed [31:0] R128_115;
wire signed [31:0] R128_138;
wire signed [31:0] R128_172;
wire signed [31:0] R128_267;
wire signed [31:0] R128_296;
wire signed [31:0] R128_416;
wire signed [31:0] R128_440;
wire signed [31:0] R129_116;
wire signed [31:0] R129_139;
wire signed [31:0] R129_173;
wire signed [31:0] R129_268;
wire signed [31:0] R129_297;
wire signed [31:0] R129_417;
wire signed [31:0] R129_441;
wire signed [31:0] R130_117;
wire signed [31:0] R130_140;
wire signed [31:0] R130_174;
wire signed [31:0] R130_269;
wire signed [31:0] R130_298;
wire signed [31:0] R130_418;
wire signed [31:0] R130_442;
wire signed [31:0] R131_118;
wire signed [31:0] R131_141;
wire signed [31:0] R131_175;
wire signed [31:0] R131_270;
wire signed [31:0] R131_299;
wire signed [31:0] R131_419;
wire signed [31:0] R131_443;
wire signed [31:0] R132_119;
wire signed [31:0] R132_142;
wire signed [31:0] R132_176;
wire signed [31:0] R132_271;
wire signed [31:0] R132_300;
wire signed [31:0] R132_420;
wire signed [31:0] R132_444;
wire signed [31:0] R133_120;
wire signed [31:0] R133_143;
wire signed [31:0] R133_177;
wire signed [31:0] R133_272;
wire signed [31:0] R133_301;
wire signed [31:0] R133_421;
wire signed [31:0] R133_445;
wire signed [31:0] R134_97;
wire signed [31:0] R134_144;
wire signed [31:0] R134_178;
wire signed [31:0] R134_273;
wire signed [31:0] R134_302;
wire signed [31:0] R134_422;
wire signed [31:0] R134_446;
wire signed [31:0] R135_98;
wire signed [31:0] R135_121;
wire signed [31:0] R135_179;
wire signed [31:0] R135_274;
wire signed [31:0] R135_303;
wire signed [31:0] R135_423;
wire signed [31:0] R135_447;
wire signed [31:0] R136_99;
wire signed [31:0] R136_122;
wire signed [31:0] R136_180;
wire signed [31:0] R136_275;
wire signed [31:0] R136_304;
wire signed [31:0] R136_424;
wire signed [31:0] R136_448;
wire signed [31:0] R137_100;
wire signed [31:0] R137_123;
wire signed [31:0] R137_181;
wire signed [31:0] R137_276;
wire signed [31:0] R137_305;
wire signed [31:0] R137_425;
wire signed [31:0] R137_449;
wire signed [31:0] R138_101;
wire signed [31:0] R138_124;
wire signed [31:0] R138_182;
wire signed [31:0] R138_277;
wire signed [31:0] R138_306;
wire signed [31:0] R138_426;
wire signed [31:0] R138_450;
wire signed [31:0] R139_102;
wire signed [31:0] R139_125;
wire signed [31:0] R139_183;
wire signed [31:0] R139_278;
wire signed [31:0] R139_307;
wire signed [31:0] R139_427;
wire signed [31:0] R139_451;
wire signed [31:0] R140_103;
wire signed [31:0] R140_126;
wire signed [31:0] R140_184;
wire signed [31:0] R140_279;
wire signed [31:0] R140_308;
wire signed [31:0] R140_428;
wire signed [31:0] R140_452;
wire signed [31:0] R141_104;
wire signed [31:0] R141_127;
wire signed [31:0] R141_185;
wire signed [31:0] R141_280;
wire signed [31:0] R141_309;
wire signed [31:0] R141_429;
wire signed [31:0] R141_453;
wire signed [31:0] R142_105;
wire signed [31:0] R142_128;
wire signed [31:0] R142_186;
wire signed [31:0] R142_281;
wire signed [31:0] R142_310;
wire signed [31:0] R142_430;
wire signed [31:0] R142_454;
wire signed [31:0] R143_106;
wire signed [31:0] R143_129;
wire signed [31:0] R143_187;
wire signed [31:0] R143_282;
wire signed [31:0] R143_311;
wire signed [31:0] R143_431;
wire signed [31:0] R143_455;
wire signed [31:0] R144_107;
wire signed [31:0] R144_130;
wire signed [31:0] R144_188;
wire signed [31:0] R144_283;
wire signed [31:0] R144_312;
wire signed [31:0] R144_432;
wire signed [31:0] R144_456;
wire signed [31:0] R145_72;
wire signed [31:0] R145_86;
wire signed [31:0] R145_220;
wire signed [31:0] R145_245;
wire signed [31:0] R145_433;
wire signed [31:0] R145_457;
wire signed [31:0] R146_49;
wire signed [31:0] R146_87;
wire signed [31:0] R146_221;
wire signed [31:0] R146_246;
wire signed [31:0] R146_434;
wire signed [31:0] R146_458;
wire signed [31:0] R147_50;
wire signed [31:0] R147_88;
wire signed [31:0] R147_222;
wire signed [31:0] R147_247;
wire signed [31:0] R147_435;
wire signed [31:0] R147_459;
wire signed [31:0] R148_51;
wire signed [31:0] R148_89;
wire signed [31:0] R148_223;
wire signed [31:0] R148_248;
wire signed [31:0] R148_436;
wire signed [31:0] R148_460;
wire signed [31:0] R149_52;
wire signed [31:0] R149_90;
wire signed [31:0] R149_224;
wire signed [31:0] R149_249;
wire signed [31:0] R149_437;
wire signed [31:0] R149_461;
wire signed [31:0] R150_53;
wire signed [31:0] R150_91;
wire signed [31:0] R150_225;
wire signed [31:0] R150_250;
wire signed [31:0] R150_438;
wire signed [31:0] R150_462;
wire signed [31:0] R151_54;
wire signed [31:0] R151_92;
wire signed [31:0] R151_226;
wire signed [31:0] R151_251;
wire signed [31:0] R151_439;
wire signed [31:0] R151_463;
wire signed [31:0] R152_55;
wire signed [31:0] R152_93;
wire signed [31:0] R152_227;
wire signed [31:0] R152_252;
wire signed [31:0] R152_440;
wire signed [31:0] R152_464;
wire signed [31:0] R153_56;
wire signed [31:0] R153_94;
wire signed [31:0] R153_228;
wire signed [31:0] R153_253;
wire signed [31:0] R153_441;
wire signed [31:0] R153_465;
wire signed [31:0] R154_57;
wire signed [31:0] R154_95;
wire signed [31:0] R154_229;
wire signed [31:0] R154_254;
wire signed [31:0] R154_442;
wire signed [31:0] R154_466;
wire signed [31:0] R155_58;
wire signed [31:0] R155_96;
wire signed [31:0] R155_230;
wire signed [31:0] R155_255;
wire signed [31:0] R155_443;
wire signed [31:0] R155_467;
wire signed [31:0] R156_59;
wire signed [31:0] R156_73;
wire signed [31:0] R156_231;
wire signed [31:0] R156_256;
wire signed [31:0] R156_444;
wire signed [31:0] R156_468;
wire signed [31:0] R157_60;
wire signed [31:0] R157_74;
wire signed [31:0] R157_232;
wire signed [31:0] R157_257;
wire signed [31:0] R157_445;
wire signed [31:0] R157_469;
wire signed [31:0] R158_61;
wire signed [31:0] R158_75;
wire signed [31:0] R158_233;
wire signed [31:0] R158_258;
wire signed [31:0] R158_446;
wire signed [31:0] R158_470;
wire signed [31:0] R159_62;
wire signed [31:0] R159_76;
wire signed [31:0] R159_234;
wire signed [31:0] R159_259;
wire signed [31:0] R159_447;
wire signed [31:0] R159_471;
wire signed [31:0] R160_63;
wire signed [31:0] R160_77;
wire signed [31:0] R160_235;
wire signed [31:0] R160_260;
wire signed [31:0] R160_448;
wire signed [31:0] R160_472;
wire signed [31:0] R161_64;
wire signed [31:0] R161_78;
wire signed [31:0] R161_236;
wire signed [31:0] R161_261;
wire signed [31:0] R161_449;
wire signed [31:0] R161_473;
wire signed [31:0] R162_65;
wire signed [31:0] R162_79;
wire signed [31:0] R162_237;
wire signed [31:0] R162_262;
wire signed [31:0] R162_450;
wire signed [31:0] R162_474;
wire signed [31:0] R163_66;
wire signed [31:0] R163_80;
wire signed [31:0] R163_238;
wire signed [31:0] R163_263;
wire signed [31:0] R163_451;
wire signed [31:0] R163_475;
wire signed [31:0] R164_67;
wire signed [31:0] R164_81;
wire signed [31:0] R164_239;
wire signed [31:0] R164_264;
wire signed [31:0] R164_452;
wire signed [31:0] R164_476;
wire signed [31:0] R165_68;
wire signed [31:0] R165_82;
wire signed [31:0] R165_240;
wire signed [31:0] R165_241;
wire signed [31:0] R165_453;
wire signed [31:0] R165_477;
wire signed [31:0] R166_69;
wire signed [31:0] R166_83;
wire signed [31:0] R166_217;
wire signed [31:0] R166_242;
wire signed [31:0] R166_454;
wire signed [31:0] R166_478;
wire signed [31:0] R167_70;
wire signed [31:0] R167_84;
wire signed [31:0] R167_218;
wire signed [31:0] R167_243;
wire signed [31:0] R167_455;
wire signed [31:0] R167_479;
wire signed [31:0] R168_71;
wire signed [31:0] R168_85;
wire signed [31:0] R168_219;
wire signed [31:0] R168_244;
wire signed [31:0] R168_456;
wire signed [31:0] R168_480;
wire signed [31:0] R169_27;
wire signed [31:0] R169_67;
wire signed [31:0] R169_145;
wire signed [31:0] R169_228;
wire signed [31:0] R169_457;
wire signed [31:0] R169_481;
wire signed [31:0] R170_28;
wire signed [31:0] R170_68;
wire signed [31:0] R170_146;
wire signed [31:0] R170_229;
wire signed [31:0] R170_458;
wire signed [31:0] R170_482;
wire signed [31:0] R171_29;
wire signed [31:0] R171_69;
wire signed [31:0] R171_147;
wire signed [31:0] R171_230;
wire signed [31:0] R171_459;
wire signed [31:0] R171_483;
wire signed [31:0] R172_30;
wire signed [31:0] R172_70;
wire signed [31:0] R172_148;
wire signed [31:0] R172_231;
wire signed [31:0] R172_460;
wire signed [31:0] R172_484;
wire signed [31:0] R173_31;
wire signed [31:0] R173_71;
wire signed [31:0] R173_149;
wire signed [31:0] R173_232;
wire signed [31:0] R173_461;
wire signed [31:0] R173_485;
wire signed [31:0] R174_32;
wire signed [31:0] R174_72;
wire signed [31:0] R174_150;
wire signed [31:0] R174_233;
wire signed [31:0] R174_462;
wire signed [31:0] R174_486;
wire signed [31:0] R175_33;
wire signed [31:0] R175_49;
wire signed [31:0] R175_151;
wire signed [31:0] R175_234;
wire signed [31:0] R175_463;
wire signed [31:0] R175_487;
wire signed [31:0] R176_34;
wire signed [31:0] R176_50;
wire signed [31:0] R176_152;
wire signed [31:0] R176_235;
wire signed [31:0] R176_464;
wire signed [31:0] R176_488;
wire signed [31:0] R177_35;
wire signed [31:0] R177_51;
wire signed [31:0] R177_153;
wire signed [31:0] R177_236;
wire signed [31:0] R177_465;
wire signed [31:0] R177_489;
wire signed [31:0] R178_36;
wire signed [31:0] R178_52;
wire signed [31:0] R178_154;
wire signed [31:0] R178_237;
wire signed [31:0] R178_466;
wire signed [31:0] R178_490;
wire signed [31:0] R179_37;
wire signed [31:0] R179_53;
wire signed [31:0] R179_155;
wire signed [31:0] R179_238;
wire signed [31:0] R179_467;
wire signed [31:0] R179_491;
wire signed [31:0] R180_38;
wire signed [31:0] R180_54;
wire signed [31:0] R180_156;
wire signed [31:0] R180_239;
wire signed [31:0] R180_468;
wire signed [31:0] R180_492;
wire signed [31:0] R181_39;
wire signed [31:0] R181_55;
wire signed [31:0] R181_157;
wire signed [31:0] R181_240;
wire signed [31:0] R181_469;
wire signed [31:0] R181_493;
wire signed [31:0] R182_40;
wire signed [31:0] R182_56;
wire signed [31:0] R182_158;
wire signed [31:0] R182_217;
wire signed [31:0] R182_470;
wire signed [31:0] R182_494;
wire signed [31:0] R183_41;
wire signed [31:0] R183_57;
wire signed [31:0] R183_159;
wire signed [31:0] R183_218;
wire signed [31:0] R183_471;
wire signed [31:0] R183_495;
wire signed [31:0] R184_42;
wire signed [31:0] R184_58;
wire signed [31:0] R184_160;
wire signed [31:0] R184_219;
wire signed [31:0] R184_472;
wire signed [31:0] R184_496;
wire signed [31:0] R185_43;
wire signed [31:0] R185_59;
wire signed [31:0] R185_161;
wire signed [31:0] R185_220;
wire signed [31:0] R185_473;
wire signed [31:0] R185_497;
wire signed [31:0] R186_44;
wire signed [31:0] R186_60;
wire signed [31:0] R186_162;
wire signed [31:0] R186_221;
wire signed [31:0] R186_474;
wire signed [31:0] R186_498;
wire signed [31:0] R187_45;
wire signed [31:0] R187_61;
wire signed [31:0] R187_163;
wire signed [31:0] R187_222;
wire signed [31:0] R187_475;
wire signed [31:0] R187_499;
wire signed [31:0] R188_46;
wire signed [31:0] R188_62;
wire signed [31:0] R188_164;
wire signed [31:0] R188_223;
wire signed [31:0] R188_476;
wire signed [31:0] R188_500;
wire signed [31:0] R189_47;
wire signed [31:0] R189_63;
wire signed [31:0] R189_165;
wire signed [31:0] R189_224;
wire signed [31:0] R189_477;
wire signed [31:0] R189_501;
wire signed [31:0] R190_48;
wire signed [31:0] R190_64;
wire signed [31:0] R190_166;
wire signed [31:0] R190_225;
wire signed [31:0] R190_478;
wire signed [31:0] R190_502;
wire signed [31:0] R191_25;
wire signed [31:0] R191_65;
wire signed [31:0] R191_167;
wire signed [31:0] R191_226;
wire signed [31:0] R191_479;
wire signed [31:0] R191_503;
wire signed [31:0] R192_26;
wire signed [31:0] R192_66;
wire signed [31:0] R192_168;
wire signed [31:0] R192_227;
wire signed [31:0] R192_480;
wire signed [31:0] R192_504;
wire signed [31:0] R193_4;
wire signed [31:0] R193_117;
wire signed [31:0] R193_127;
wire signed [31:0] R193_179;
wire signed [31:0] R193_277;
wire signed [31:0] R193_481;
wire signed [31:0] R193_505;
wire signed [31:0] R194_5;
wire signed [31:0] R194_118;
wire signed [31:0] R194_128;
wire signed [31:0] R194_180;
wire signed [31:0] R194_278;
wire signed [31:0] R194_482;
wire signed [31:0] R194_506;
wire signed [31:0] R195_6;
wire signed [31:0] R195_119;
wire signed [31:0] R195_129;
wire signed [31:0] R195_181;
wire signed [31:0] R195_279;
wire signed [31:0] R195_483;
wire signed [31:0] R195_507;
wire signed [31:0] R196_7;
wire signed [31:0] R196_120;
wire signed [31:0] R196_130;
wire signed [31:0] R196_182;
wire signed [31:0] R196_280;
wire signed [31:0] R196_484;
wire signed [31:0] R196_508;
wire signed [31:0] R197_8;
wire signed [31:0] R197_97;
wire signed [31:0] R197_131;
wire signed [31:0] R197_183;
wire signed [31:0] R197_281;
wire signed [31:0] R197_485;
wire signed [31:0] R197_509;
wire signed [31:0] R198_9;
wire signed [31:0] R198_98;
wire signed [31:0] R198_132;
wire signed [31:0] R198_184;
wire signed [31:0] R198_282;
wire signed [31:0] R198_486;
wire signed [31:0] R198_510;
wire signed [31:0] R199_10;
wire signed [31:0] R199_99;
wire signed [31:0] R199_133;
wire signed [31:0] R199_185;
wire signed [31:0] R199_283;
wire signed [31:0] R199_487;
wire signed [31:0] R199_511;
wire signed [31:0] R200_11;
wire signed [31:0] R200_100;
wire signed [31:0] R200_134;
wire signed [31:0] R200_186;
wire signed [31:0] R200_284;
wire signed [31:0] R200_488;
wire signed [31:0] R200_512;
wire signed [31:0] R201_12;
wire signed [31:0] R201_101;
wire signed [31:0] R201_135;
wire signed [31:0] R201_187;
wire signed [31:0] R201_285;
wire signed [31:0] R201_489;
wire signed [31:0] R201_513;
wire signed [31:0] R202_13;
wire signed [31:0] R202_102;
wire signed [31:0] R202_136;
wire signed [31:0] R202_188;
wire signed [31:0] R202_286;
wire signed [31:0] R202_490;
wire signed [31:0] R202_514;
wire signed [31:0] R203_14;
wire signed [31:0] R203_103;
wire signed [31:0] R203_137;
wire signed [31:0] R203_189;
wire signed [31:0] R203_287;
wire signed [31:0] R203_491;
wire signed [31:0] R203_515;
wire signed [31:0] R204_15;
wire signed [31:0] R204_104;
wire signed [31:0] R204_138;
wire signed [31:0] R204_190;
wire signed [31:0] R204_288;
wire signed [31:0] R204_492;
wire signed [31:0] R204_516;
wire signed [31:0] R205_16;
wire signed [31:0] R205_105;
wire signed [31:0] R205_139;
wire signed [31:0] R205_191;
wire signed [31:0] R205_265;
wire signed [31:0] R205_493;
wire signed [31:0] R205_517;
wire signed [31:0] R206_17;
wire signed [31:0] R206_106;
wire signed [31:0] R206_140;
wire signed [31:0] R206_192;
wire signed [31:0] R206_266;
wire signed [31:0] R206_494;
wire signed [31:0] R206_518;
wire signed [31:0] R207_18;
wire signed [31:0] R207_107;
wire signed [31:0] R207_141;
wire signed [31:0] R207_169;
wire signed [31:0] R207_267;
wire signed [31:0] R207_495;
wire signed [31:0] R207_519;
wire signed [31:0] R208_19;
wire signed [31:0] R208_108;
wire signed [31:0] R208_142;
wire signed [31:0] R208_170;
wire signed [31:0] R208_268;
wire signed [31:0] R208_496;
wire signed [31:0] R208_520;
wire signed [31:0] R209_20;
wire signed [31:0] R209_109;
wire signed [31:0] R209_143;
wire signed [31:0] R209_171;
wire signed [31:0] R209_269;
wire signed [31:0] R209_497;
wire signed [31:0] R209_521;
wire signed [31:0] R210_21;
wire signed [31:0] R210_110;
wire signed [31:0] R210_144;
wire signed [31:0] R210_172;
wire signed [31:0] R210_270;
wire signed [31:0] R210_498;
wire signed [31:0] R210_522;
wire signed [31:0] R211_22;
wire signed [31:0] R211_111;
wire signed [31:0] R211_121;
wire signed [31:0] R211_173;
wire signed [31:0] R211_271;
wire signed [31:0] R211_499;
wire signed [31:0] R211_523;
wire signed [31:0] R212_23;
wire signed [31:0] R212_112;
wire signed [31:0] R212_122;
wire signed [31:0] R212_174;
wire signed [31:0] R212_272;
wire signed [31:0] R212_500;
wire signed [31:0] R212_524;
wire signed [31:0] R213_24;
wire signed [31:0] R213_113;
wire signed [31:0] R213_123;
wire signed [31:0] R213_175;
wire signed [31:0] R213_273;
wire signed [31:0] R213_501;
wire signed [31:0] R213_525;
wire signed [31:0] R214_1;
wire signed [31:0] R214_114;
wire signed [31:0] R214_124;
wire signed [31:0] R214_176;
wire signed [31:0] R214_274;
wire signed [31:0] R214_502;
wire signed [31:0] R214_526;
wire signed [31:0] R215_2;
wire signed [31:0] R215_115;
wire signed [31:0] R215_125;
wire signed [31:0] R215_177;
wire signed [31:0] R215_275;
wire signed [31:0] R215_503;
wire signed [31:0] R215_527;
wire signed [31:0] R216_3;
wire signed [31:0] R216_116;
wire signed [31:0] R216_126;
wire signed [31:0] R216_178;
wire signed [31:0] R216_276;
wire signed [31:0] R216_504;
wire signed [31:0] R216_528;
wire signed [31:0] R217_144;
wire signed [31:0] R217_183;
wire signed [31:0] R217_258;
wire signed [31:0] R217_283;
wire signed [31:0] R217_505;
wire signed [31:0] R217_529;
wire signed [31:0] R218_121;
wire signed [31:0] R218_184;
wire signed [31:0] R218_259;
wire signed [31:0] R218_284;
wire signed [31:0] R218_506;
wire signed [31:0] R218_530;
wire signed [31:0] R219_122;
wire signed [31:0] R219_185;
wire signed [31:0] R219_260;
wire signed [31:0] R219_285;
wire signed [31:0] R219_507;
wire signed [31:0] R219_531;
wire signed [31:0] R220_123;
wire signed [31:0] R220_186;
wire signed [31:0] R220_261;
wire signed [31:0] R220_286;
wire signed [31:0] R220_508;
wire signed [31:0] R220_532;
wire signed [31:0] R221_124;
wire signed [31:0] R221_187;
wire signed [31:0] R221_262;
wire signed [31:0] R221_287;
wire signed [31:0] R221_509;
wire signed [31:0] R221_533;
wire signed [31:0] R222_125;
wire signed [31:0] R222_188;
wire signed [31:0] R222_263;
wire signed [31:0] R222_288;
wire signed [31:0] R222_510;
wire signed [31:0] R222_534;
wire signed [31:0] R223_126;
wire signed [31:0] R223_189;
wire signed [31:0] R223_264;
wire signed [31:0] R223_265;
wire signed [31:0] R223_511;
wire signed [31:0] R223_535;
wire signed [31:0] R224_127;
wire signed [31:0] R224_190;
wire signed [31:0] R224_241;
wire signed [31:0] R224_266;
wire signed [31:0] R224_512;
wire signed [31:0] R224_536;
wire signed [31:0] R225_128;
wire signed [31:0] R225_191;
wire signed [31:0] R225_242;
wire signed [31:0] R225_267;
wire signed [31:0] R225_513;
wire signed [31:0] R225_537;
wire signed [31:0] R226_129;
wire signed [31:0] R226_192;
wire signed [31:0] R226_243;
wire signed [31:0] R226_268;
wire signed [31:0] R226_514;
wire signed [31:0] R226_538;
wire signed [31:0] R227_130;
wire signed [31:0] R227_169;
wire signed [31:0] R227_244;
wire signed [31:0] R227_269;
wire signed [31:0] R227_515;
wire signed [31:0] R227_539;
wire signed [31:0] R228_131;
wire signed [31:0] R228_170;
wire signed [31:0] R228_245;
wire signed [31:0] R228_270;
wire signed [31:0] R228_516;
wire signed [31:0] R228_540;
wire signed [31:0] R229_132;
wire signed [31:0] R229_171;
wire signed [31:0] R229_246;
wire signed [31:0] R229_271;
wire signed [31:0] R229_517;
wire signed [31:0] R229_541;
wire signed [31:0] R230_133;
wire signed [31:0] R230_172;
wire signed [31:0] R230_247;
wire signed [31:0] R230_272;
wire signed [31:0] R230_518;
wire signed [31:0] R230_542;
wire signed [31:0] R231_134;
wire signed [31:0] R231_173;
wire signed [31:0] R231_248;
wire signed [31:0] R231_273;
wire signed [31:0] R231_519;
wire signed [31:0] R231_543;
wire signed [31:0] R232_135;
wire signed [31:0] R232_174;
wire signed [31:0] R232_249;
wire signed [31:0] R232_274;
wire signed [31:0] R232_520;
wire signed [31:0] R232_544;
wire signed [31:0] R233_136;
wire signed [31:0] R233_175;
wire signed [31:0] R233_250;
wire signed [31:0] R233_275;
wire signed [31:0] R233_521;
wire signed [31:0] R233_545;
wire signed [31:0] R234_137;
wire signed [31:0] R234_176;
wire signed [31:0] R234_251;
wire signed [31:0] R234_276;
wire signed [31:0] R234_522;
wire signed [31:0] R234_546;
wire signed [31:0] R235_138;
wire signed [31:0] R235_177;
wire signed [31:0] R235_252;
wire signed [31:0] R235_277;
wire signed [31:0] R235_523;
wire signed [31:0] R235_547;
wire signed [31:0] R236_139;
wire signed [31:0] R236_178;
wire signed [31:0] R236_253;
wire signed [31:0] R236_278;
wire signed [31:0] R236_524;
wire signed [31:0] R236_548;
wire signed [31:0] R237_140;
wire signed [31:0] R237_179;
wire signed [31:0] R237_254;
wire signed [31:0] R237_279;
wire signed [31:0] R237_525;
wire signed [31:0] R237_549;
wire signed [31:0] R238_141;
wire signed [31:0] R238_180;
wire signed [31:0] R238_255;
wire signed [31:0] R238_280;
wire signed [31:0] R238_526;
wire signed [31:0] R238_550;
wire signed [31:0] R239_142;
wire signed [31:0] R239_181;
wire signed [31:0] R239_256;
wire signed [31:0] R239_281;
wire signed [31:0] R239_527;
wire signed [31:0] R239_551;
wire signed [31:0] R240_143;
wire signed [31:0] R240_182;
wire signed [31:0] R240_257;
wire signed [31:0] R240_282;
wire signed [31:0] R240_528;
wire signed [31:0] R240_552;
wire signed [31:0] R241_50;
wire signed [31:0] R241_89;
wire signed [31:0] R241_202;
wire signed [31:0] R241_229;
wire signed [31:0] R241_529;
wire signed [31:0] R241_553;
wire signed [31:0] R242_51;
wire signed [31:0] R242_90;
wire signed [31:0] R242_203;
wire signed [31:0] R242_230;
wire signed [31:0] R242_530;
wire signed [31:0] R242_554;
wire signed [31:0] R243_52;
wire signed [31:0] R243_91;
wire signed [31:0] R243_204;
wire signed [31:0] R243_231;
wire signed [31:0] R243_531;
wire signed [31:0] R243_555;
wire signed [31:0] R244_53;
wire signed [31:0] R244_92;
wire signed [31:0] R244_205;
wire signed [31:0] R244_232;
wire signed [31:0] R244_532;
wire signed [31:0] R244_556;
wire signed [31:0] R245_54;
wire signed [31:0] R245_93;
wire signed [31:0] R245_206;
wire signed [31:0] R245_233;
wire signed [31:0] R245_533;
wire signed [31:0] R245_557;
wire signed [31:0] R246_55;
wire signed [31:0] R246_94;
wire signed [31:0] R246_207;
wire signed [31:0] R246_234;
wire signed [31:0] R246_534;
wire signed [31:0] R246_558;
wire signed [31:0] R247_56;
wire signed [31:0] R247_95;
wire signed [31:0] R247_208;
wire signed [31:0] R247_235;
wire signed [31:0] R247_535;
wire signed [31:0] R247_559;
wire signed [31:0] R248_57;
wire signed [31:0] R248_96;
wire signed [31:0] R248_209;
wire signed [31:0] R248_236;
wire signed [31:0] R248_536;
wire signed [31:0] R248_560;
wire signed [31:0] R249_58;
wire signed [31:0] R249_73;
wire signed [31:0] R249_210;
wire signed [31:0] R249_237;
wire signed [31:0] R249_537;
wire signed [31:0] R249_561;
wire signed [31:0] R250_59;
wire signed [31:0] R250_74;
wire signed [31:0] R250_211;
wire signed [31:0] R250_238;
wire signed [31:0] R250_538;
wire signed [31:0] R250_562;
wire signed [31:0] R251_60;
wire signed [31:0] R251_75;
wire signed [31:0] R251_212;
wire signed [31:0] R251_239;
wire signed [31:0] R251_539;
wire signed [31:0] R251_563;
wire signed [31:0] R252_61;
wire signed [31:0] R252_76;
wire signed [31:0] R252_213;
wire signed [31:0] R252_240;
wire signed [31:0] R252_540;
wire signed [31:0] R252_564;
wire signed [31:0] R253_62;
wire signed [31:0] R253_77;
wire signed [31:0] R253_214;
wire signed [31:0] R253_217;
wire signed [31:0] R253_541;
wire signed [31:0] R253_565;
wire signed [31:0] R254_63;
wire signed [31:0] R254_78;
wire signed [31:0] R254_215;
wire signed [31:0] R254_218;
wire signed [31:0] R254_542;
wire signed [31:0] R254_566;
wire signed [31:0] R255_64;
wire signed [31:0] R255_79;
wire signed [31:0] R255_216;
wire signed [31:0] R255_219;
wire signed [31:0] R255_543;
wire signed [31:0] R255_567;
wire signed [31:0] R256_65;
wire signed [31:0] R256_80;
wire signed [31:0] R256_193;
wire signed [31:0] R256_220;
wire signed [31:0] R256_544;
wire signed [31:0] R256_568;
wire signed [31:0] R257_66;
wire signed [31:0] R257_81;
wire signed [31:0] R257_194;
wire signed [31:0] R257_221;
wire signed [31:0] R257_545;
wire signed [31:0] R257_569;
wire signed [31:0] R258_67;
wire signed [31:0] R258_82;
wire signed [31:0] R258_195;
wire signed [31:0] R258_222;
wire signed [31:0] R258_546;
wire signed [31:0] R258_570;
wire signed [31:0] R259_68;
wire signed [31:0] R259_83;
wire signed [31:0] R259_196;
wire signed [31:0] R259_223;
wire signed [31:0] R259_547;
wire signed [31:0] R259_571;
wire signed [31:0] R260_69;
wire signed [31:0] R260_84;
wire signed [31:0] R260_197;
wire signed [31:0] R260_224;
wire signed [31:0] R260_548;
wire signed [31:0] R260_572;
wire signed [31:0] R261_70;
wire signed [31:0] R261_85;
wire signed [31:0] R261_198;
wire signed [31:0] R261_225;
wire signed [31:0] R261_549;
wire signed [31:0] R261_573;
wire signed [31:0] R262_71;
wire signed [31:0] R262_86;
wire signed [31:0] R262_199;
wire signed [31:0] R262_226;
wire signed [31:0] R262_550;
wire signed [31:0] R262_574;
wire signed [31:0] R263_72;
wire signed [31:0] R263_87;
wire signed [31:0] R263_200;
wire signed [31:0] R263_227;
wire signed [31:0] R263_551;
wire signed [31:0] R263_575;
wire signed [31:0] R264_49;
wire signed [31:0] R264_88;
wire signed [31:0] R264_201;
wire signed [31:0] R264_228;
wire signed [31:0] R264_552;
wire signed [31:0] R264_576;
wire signed [31:0] R265_11;
wire signed [31:0] R265_137;
wire signed [31:0] R265_179;
wire signed [31:0] R265_271;
wire signed [31:0] R265_290;
wire signed [31:0] R265_553;
wire signed [31:0] R266_12;
wire signed [31:0] R266_138;
wire signed [31:0] R266_180;
wire signed [31:0] R266_272;
wire signed [31:0] R266_291;
wire signed [31:0] R266_554;
wire signed [31:0] R267_13;
wire signed [31:0] R267_139;
wire signed [31:0] R267_181;
wire signed [31:0] R267_273;
wire signed [31:0] R267_292;
wire signed [31:0] R267_555;
wire signed [31:0] R268_14;
wire signed [31:0] R268_140;
wire signed [31:0] R268_182;
wire signed [31:0] R268_274;
wire signed [31:0] R268_293;
wire signed [31:0] R268_556;
wire signed [31:0] R269_15;
wire signed [31:0] R269_141;
wire signed [31:0] R269_183;
wire signed [31:0] R269_275;
wire signed [31:0] R269_294;
wire signed [31:0] R269_557;
wire signed [31:0] R270_16;
wire signed [31:0] R270_142;
wire signed [31:0] R270_184;
wire signed [31:0] R270_276;
wire signed [31:0] R270_295;
wire signed [31:0] R270_558;
wire signed [31:0] R271_17;
wire signed [31:0] R271_143;
wire signed [31:0] R271_185;
wire signed [31:0] R271_277;
wire signed [31:0] R271_296;
wire signed [31:0] R271_559;
wire signed [31:0] R272_18;
wire signed [31:0] R272_144;
wire signed [31:0] R272_186;
wire signed [31:0] R272_278;
wire signed [31:0] R272_297;
wire signed [31:0] R272_560;
wire signed [31:0] R273_19;
wire signed [31:0] R273_121;
wire signed [31:0] R273_187;
wire signed [31:0] R273_279;
wire signed [31:0] R273_298;
wire signed [31:0] R273_561;
wire signed [31:0] R274_20;
wire signed [31:0] R274_122;
wire signed [31:0] R274_188;
wire signed [31:0] R274_280;
wire signed [31:0] R274_299;
wire signed [31:0] R274_562;
wire signed [31:0] R275_21;
wire signed [31:0] R275_123;
wire signed [31:0] R275_189;
wire signed [31:0] R275_281;
wire signed [31:0] R275_300;
wire signed [31:0] R275_563;
wire signed [31:0] R276_22;
wire signed [31:0] R276_124;
wire signed [31:0] R276_190;
wire signed [31:0] R276_282;
wire signed [31:0] R276_301;
wire signed [31:0] R276_564;
wire signed [31:0] R277_23;
wire signed [31:0] R277_125;
wire signed [31:0] R277_191;
wire signed [31:0] R277_283;
wire signed [31:0] R277_302;
wire signed [31:0] R277_565;
wire signed [31:0] R278_24;
wire signed [31:0] R278_126;
wire signed [31:0] R278_192;
wire signed [31:0] R278_284;
wire signed [31:0] R278_303;
wire signed [31:0] R278_566;
wire signed [31:0] R279_1;
wire signed [31:0] R279_127;
wire signed [31:0] R279_169;
wire signed [31:0] R279_285;
wire signed [31:0] R279_304;
wire signed [31:0] R279_567;
wire signed [31:0] R280_2;
wire signed [31:0] R280_128;
wire signed [31:0] R280_170;
wire signed [31:0] R280_286;
wire signed [31:0] R280_305;
wire signed [31:0] R280_568;
wire signed [31:0] R281_3;
wire signed [31:0] R281_129;
wire signed [31:0] R281_171;
wire signed [31:0] R281_287;
wire signed [31:0] R281_306;
wire signed [31:0] R281_569;
wire signed [31:0] R282_4;
wire signed [31:0] R282_130;
wire signed [31:0] R282_172;
wire signed [31:0] R282_288;
wire signed [31:0] R282_307;
wire signed [31:0] R282_570;
wire signed [31:0] R283_5;
wire signed [31:0] R283_131;
wire signed [31:0] R283_173;
wire signed [31:0] R283_265;
wire signed [31:0] R283_308;
wire signed [31:0] R283_571;
wire signed [31:0] R284_6;
wire signed [31:0] R284_132;
wire signed [31:0] R284_174;
wire signed [31:0] R284_266;
wire signed [31:0] R284_309;
wire signed [31:0] R284_572;
wire signed [31:0] R285_7;
wire signed [31:0] R285_133;
wire signed [31:0] R285_175;
wire signed [31:0] R285_267;
wire signed [31:0] R285_310;
wire signed [31:0] R285_573;
wire signed [31:0] R286_8;
wire signed [31:0] R286_134;
wire signed [31:0] R286_176;
wire signed [31:0] R286_268;
wire signed [31:0] R286_311;
wire signed [31:0] R286_574;
wire signed [31:0] R287_9;
wire signed [31:0] R287_135;
wire signed [31:0] R287_177;
wire signed [31:0] R287_269;
wire signed [31:0] R287_312;
wire signed [31:0] R287_575;
wire signed [31:0] R288_10;
wire signed [31:0] R288_136;
wire signed [31:0] R288_178;
wire signed [31:0] R288_270;
wire signed [31:0] R288_289;
wire signed [31:0] R288_576;
wire signed [31:0] Q1_48;
wire signed [31:0] Q1_67;
wire signed [31:0] Q1_206;
wire signed [31:0] Q1_237;
wire signed [31:0] Q1_290;
wire signed [31:0] Q1_313;
wire signed [31:0] Q2_25;
wire signed [31:0] Q2_68;
wire signed [31:0] Q2_207;
wire signed [31:0] Q2_238;
wire signed [31:0] Q2_291;
wire signed [31:0] Q2_314;
wire signed [31:0] Q3_26;
wire signed [31:0] Q3_69;
wire signed [31:0] Q3_208;
wire signed [31:0] Q3_239;
wire signed [31:0] Q3_292;
wire signed [31:0] Q3_315;
wire signed [31:0] Q4_27;
wire signed [31:0] Q4_70;
wire signed [31:0] Q4_209;
wire signed [31:0] Q4_240;
wire signed [31:0] Q4_293;
wire signed [31:0] Q4_316;
wire signed [31:0] Q5_28;
wire signed [31:0] Q5_71;
wire signed [31:0] Q5_210;
wire signed [31:0] Q5_217;
wire signed [31:0] Q5_294;
wire signed [31:0] Q5_317;
wire signed [31:0] Q6_29;
wire signed [31:0] Q6_72;
wire signed [31:0] Q6_211;
wire signed [31:0] Q6_218;
wire signed [31:0] Q6_295;
wire signed [31:0] Q6_318;
wire signed [31:0] Q7_30;
wire signed [31:0] Q7_49;
wire signed [31:0] Q7_212;
wire signed [31:0] Q7_219;
wire signed [31:0] Q7_296;
wire signed [31:0] Q7_319;
wire signed [31:0] Q8_31;
wire signed [31:0] Q8_50;
wire signed [31:0] Q8_213;
wire signed [31:0] Q8_220;
wire signed [31:0] Q8_297;
wire signed [31:0] Q8_320;
wire signed [31:0] Q9_32;
wire signed [31:0] Q9_51;
wire signed [31:0] Q9_214;
wire signed [31:0] Q9_221;
wire signed [31:0] Q9_298;
wire signed [31:0] Q9_321;
wire signed [31:0] Q10_33;
wire signed [31:0] Q10_52;
wire signed [31:0] Q10_215;
wire signed [31:0] Q10_222;
wire signed [31:0] Q10_299;
wire signed [31:0] Q10_322;
wire signed [31:0] Q11_34;
wire signed [31:0] Q11_53;
wire signed [31:0] Q11_216;
wire signed [31:0] Q11_223;
wire signed [31:0] Q11_300;
wire signed [31:0] Q11_323;
wire signed [31:0] Q12_35;
wire signed [31:0] Q12_54;
wire signed [31:0] Q12_193;
wire signed [31:0] Q12_224;
wire signed [31:0] Q12_301;
wire signed [31:0] Q12_324;
wire signed [31:0] Q13_36;
wire signed [31:0] Q13_55;
wire signed [31:0] Q13_194;
wire signed [31:0] Q13_225;
wire signed [31:0] Q13_302;
wire signed [31:0] Q13_325;
wire signed [31:0] Q14_37;
wire signed [31:0] Q14_56;
wire signed [31:0] Q14_195;
wire signed [31:0] Q14_226;
wire signed [31:0] Q14_303;
wire signed [31:0] Q14_326;
wire signed [31:0] Q15_38;
wire signed [31:0] Q15_57;
wire signed [31:0] Q15_196;
wire signed [31:0] Q15_227;
wire signed [31:0] Q15_304;
wire signed [31:0] Q15_327;
wire signed [31:0] Q16_39;
wire signed [31:0] Q16_58;
wire signed [31:0] Q16_197;
wire signed [31:0] Q16_228;
wire signed [31:0] Q16_305;
wire signed [31:0] Q16_328;
wire signed [31:0] Q17_40;
wire signed [31:0] Q17_59;
wire signed [31:0] Q17_198;
wire signed [31:0] Q17_229;
wire signed [31:0] Q17_306;
wire signed [31:0] Q17_329;
wire signed [31:0] Q18_41;
wire signed [31:0] Q18_60;
wire signed [31:0] Q18_199;
wire signed [31:0] Q18_230;
wire signed [31:0] Q18_307;
wire signed [31:0] Q18_330;
wire signed [31:0] Q19_42;
wire signed [31:0] Q19_61;
wire signed [31:0] Q19_200;
wire signed [31:0] Q19_231;
wire signed [31:0] Q19_308;
wire signed [31:0] Q19_331;
wire signed [31:0] Q20_43;
wire signed [31:0] Q20_62;
wire signed [31:0] Q20_201;
wire signed [31:0] Q20_232;
wire signed [31:0] Q20_309;
wire signed [31:0] Q20_332;
wire signed [31:0] Q21_44;
wire signed [31:0] Q21_63;
wire signed [31:0] Q21_202;
wire signed [31:0] Q21_233;
wire signed [31:0] Q21_310;
wire signed [31:0] Q21_333;
wire signed [31:0] Q22_45;
wire signed [31:0] Q22_64;
wire signed [31:0] Q22_203;
wire signed [31:0] Q22_234;
wire signed [31:0] Q22_311;
wire signed [31:0] Q22_334;
wire signed [31:0] Q23_46;
wire signed [31:0] Q23_65;
wire signed [31:0] Q23_204;
wire signed [31:0] Q23_235;
wire signed [31:0] Q23_312;
wire signed [31:0] Q23_335;
wire signed [31:0] Q24_47;
wire signed [31:0] Q24_66;
wire signed [31:0] Q24_205;
wire signed [31:0] Q24_236;
wire signed [31:0] Q24_289;
wire signed [31:0] Q24_336;
wire signed [31:0] Q25_31;
wire signed [31:0] Q25_126;
wire signed [31:0] Q25_164;
wire signed [31:0] Q25_171;
wire signed [31:0] Q25_268;
wire signed [31:0] Q25_313;
wire signed [31:0] Q25_337;
wire signed [31:0] Q26_32;
wire signed [31:0] Q26_127;
wire signed [31:0] Q26_165;
wire signed [31:0] Q26_172;
wire signed [31:0] Q26_269;
wire signed [31:0] Q26_314;
wire signed [31:0] Q26_338;
wire signed [31:0] Q27_33;
wire signed [31:0] Q27_128;
wire signed [31:0] Q27_166;
wire signed [31:0] Q27_173;
wire signed [31:0] Q27_270;
wire signed [31:0] Q27_315;
wire signed [31:0] Q27_339;
wire signed [31:0] Q28_34;
wire signed [31:0] Q28_129;
wire signed [31:0] Q28_167;
wire signed [31:0] Q28_174;
wire signed [31:0] Q28_271;
wire signed [31:0] Q28_316;
wire signed [31:0] Q28_340;
wire signed [31:0] Q29_35;
wire signed [31:0] Q29_130;
wire signed [31:0] Q29_168;
wire signed [31:0] Q29_175;
wire signed [31:0] Q29_272;
wire signed [31:0] Q29_317;
wire signed [31:0] Q29_341;
wire signed [31:0] Q30_36;
wire signed [31:0] Q30_131;
wire signed [31:0] Q30_145;
wire signed [31:0] Q30_176;
wire signed [31:0] Q30_273;
wire signed [31:0] Q30_318;
wire signed [31:0] Q30_342;
wire signed [31:0] Q31_37;
wire signed [31:0] Q31_132;
wire signed [31:0] Q31_146;
wire signed [31:0] Q31_177;
wire signed [31:0] Q31_274;
wire signed [31:0] Q31_319;
wire signed [31:0] Q31_343;
wire signed [31:0] Q32_38;
wire signed [31:0] Q32_133;
wire signed [31:0] Q32_147;
wire signed [31:0] Q32_178;
wire signed [31:0] Q32_275;
wire signed [31:0] Q32_320;
wire signed [31:0] Q32_344;
wire signed [31:0] Q33_39;
wire signed [31:0] Q33_134;
wire signed [31:0] Q33_148;
wire signed [31:0] Q33_179;
wire signed [31:0] Q33_276;
wire signed [31:0] Q33_321;
wire signed [31:0] Q33_345;
wire signed [31:0] Q34_40;
wire signed [31:0] Q34_135;
wire signed [31:0] Q34_149;
wire signed [31:0] Q34_180;
wire signed [31:0] Q34_277;
wire signed [31:0] Q34_322;
wire signed [31:0] Q34_346;
wire signed [31:0] Q35_41;
wire signed [31:0] Q35_136;
wire signed [31:0] Q35_150;
wire signed [31:0] Q35_181;
wire signed [31:0] Q35_278;
wire signed [31:0] Q35_323;
wire signed [31:0] Q35_347;
wire signed [31:0] Q36_42;
wire signed [31:0] Q36_137;
wire signed [31:0] Q36_151;
wire signed [31:0] Q36_182;
wire signed [31:0] Q36_279;
wire signed [31:0] Q36_324;
wire signed [31:0] Q36_348;
wire signed [31:0] Q37_43;
wire signed [31:0] Q37_138;
wire signed [31:0] Q37_152;
wire signed [31:0] Q37_183;
wire signed [31:0] Q37_280;
wire signed [31:0] Q37_325;
wire signed [31:0] Q37_349;
wire signed [31:0] Q38_44;
wire signed [31:0] Q38_139;
wire signed [31:0] Q38_153;
wire signed [31:0] Q38_184;
wire signed [31:0] Q38_281;
wire signed [31:0] Q38_326;
wire signed [31:0] Q38_350;
wire signed [31:0] Q39_45;
wire signed [31:0] Q39_140;
wire signed [31:0] Q39_154;
wire signed [31:0] Q39_185;
wire signed [31:0] Q39_282;
wire signed [31:0] Q39_327;
wire signed [31:0] Q39_351;
wire signed [31:0] Q40_46;
wire signed [31:0] Q40_141;
wire signed [31:0] Q40_155;
wire signed [31:0] Q40_186;
wire signed [31:0] Q40_283;
wire signed [31:0] Q40_328;
wire signed [31:0] Q40_352;
wire signed [31:0] Q41_47;
wire signed [31:0] Q41_142;
wire signed [31:0] Q41_156;
wire signed [31:0] Q41_187;
wire signed [31:0] Q41_284;
wire signed [31:0] Q41_329;
wire signed [31:0] Q41_353;
wire signed [31:0] Q42_48;
wire signed [31:0] Q42_143;
wire signed [31:0] Q42_157;
wire signed [31:0] Q42_188;
wire signed [31:0] Q42_285;
wire signed [31:0] Q42_330;
wire signed [31:0] Q42_354;
wire signed [31:0] Q43_25;
wire signed [31:0] Q43_144;
wire signed [31:0] Q43_158;
wire signed [31:0] Q43_189;
wire signed [31:0] Q43_286;
wire signed [31:0] Q43_331;
wire signed [31:0] Q43_355;
wire signed [31:0] Q44_26;
wire signed [31:0] Q44_121;
wire signed [31:0] Q44_159;
wire signed [31:0] Q44_190;
wire signed [31:0] Q44_287;
wire signed [31:0] Q44_332;
wire signed [31:0] Q44_356;
wire signed [31:0] Q45_27;
wire signed [31:0] Q45_122;
wire signed [31:0] Q45_160;
wire signed [31:0] Q45_191;
wire signed [31:0] Q45_288;
wire signed [31:0] Q45_333;
wire signed [31:0] Q45_357;
wire signed [31:0] Q46_28;
wire signed [31:0] Q46_123;
wire signed [31:0] Q46_161;
wire signed [31:0] Q46_192;
wire signed [31:0] Q46_265;
wire signed [31:0] Q46_334;
wire signed [31:0] Q46_358;
wire signed [31:0] Q47_29;
wire signed [31:0] Q47_124;
wire signed [31:0] Q47_162;
wire signed [31:0] Q47_169;
wire signed [31:0] Q47_266;
wire signed [31:0] Q47_335;
wire signed [31:0] Q47_359;
wire signed [31:0] Q48_30;
wire signed [31:0] Q48_125;
wire signed [31:0] Q48_163;
wire signed [31:0] Q48_170;
wire signed [31:0] Q48_267;
wire signed [31:0] Q48_336;
wire signed [31:0] Q48_360;
wire signed [31:0] Q49_79;
wire signed [31:0] Q49_102;
wire signed [31:0] Q49_141;
wire signed [31:0] Q49_177;
wire signed [31:0] Q49_265;
wire signed [31:0] Q49_337;
wire signed [31:0] Q49_361;
wire signed [31:0] Q50_80;
wire signed [31:0] Q50_103;
wire signed [31:0] Q50_142;
wire signed [31:0] Q50_178;
wire signed [31:0] Q50_266;
wire signed [31:0] Q50_338;
wire signed [31:0] Q50_362;
wire signed [31:0] Q51_81;
wire signed [31:0] Q51_104;
wire signed [31:0] Q51_143;
wire signed [31:0] Q51_179;
wire signed [31:0] Q51_267;
wire signed [31:0] Q51_339;
wire signed [31:0] Q51_363;
wire signed [31:0] Q52_82;
wire signed [31:0] Q52_105;
wire signed [31:0] Q52_144;
wire signed [31:0] Q52_180;
wire signed [31:0] Q52_268;
wire signed [31:0] Q52_340;
wire signed [31:0] Q52_364;
wire signed [31:0] Q53_83;
wire signed [31:0] Q53_106;
wire signed [31:0] Q53_121;
wire signed [31:0] Q53_181;
wire signed [31:0] Q53_269;
wire signed [31:0] Q53_341;
wire signed [31:0] Q53_365;
wire signed [31:0] Q54_84;
wire signed [31:0] Q54_107;
wire signed [31:0] Q54_122;
wire signed [31:0] Q54_182;
wire signed [31:0] Q54_270;
wire signed [31:0] Q54_342;
wire signed [31:0] Q54_366;
wire signed [31:0] Q55_85;
wire signed [31:0] Q55_108;
wire signed [31:0] Q55_123;
wire signed [31:0] Q55_183;
wire signed [31:0] Q55_271;
wire signed [31:0] Q55_343;
wire signed [31:0] Q55_367;
wire signed [31:0] Q56_86;
wire signed [31:0] Q56_109;
wire signed [31:0] Q56_124;
wire signed [31:0] Q56_184;
wire signed [31:0] Q56_272;
wire signed [31:0] Q56_344;
wire signed [31:0] Q56_368;
wire signed [31:0] Q57_87;
wire signed [31:0] Q57_110;
wire signed [31:0] Q57_125;
wire signed [31:0] Q57_185;
wire signed [31:0] Q57_273;
wire signed [31:0] Q57_345;
wire signed [31:0] Q57_369;
wire signed [31:0] Q58_88;
wire signed [31:0] Q58_111;
wire signed [31:0] Q58_126;
wire signed [31:0] Q58_186;
wire signed [31:0] Q58_274;
wire signed [31:0] Q58_346;
wire signed [31:0] Q58_370;
wire signed [31:0] Q59_89;
wire signed [31:0] Q59_112;
wire signed [31:0] Q59_127;
wire signed [31:0] Q59_187;
wire signed [31:0] Q59_275;
wire signed [31:0] Q59_347;
wire signed [31:0] Q59_371;
wire signed [31:0] Q60_90;
wire signed [31:0] Q60_113;
wire signed [31:0] Q60_128;
wire signed [31:0] Q60_188;
wire signed [31:0] Q60_276;
wire signed [31:0] Q60_348;
wire signed [31:0] Q60_372;
wire signed [31:0] Q61_91;
wire signed [31:0] Q61_114;
wire signed [31:0] Q61_129;
wire signed [31:0] Q61_189;
wire signed [31:0] Q61_277;
wire signed [31:0] Q61_349;
wire signed [31:0] Q61_373;
wire signed [31:0] Q62_92;
wire signed [31:0] Q62_115;
wire signed [31:0] Q62_130;
wire signed [31:0] Q62_190;
wire signed [31:0] Q62_278;
wire signed [31:0] Q62_350;
wire signed [31:0] Q62_374;
wire signed [31:0] Q63_93;
wire signed [31:0] Q63_116;
wire signed [31:0] Q63_131;
wire signed [31:0] Q63_191;
wire signed [31:0] Q63_279;
wire signed [31:0] Q63_351;
wire signed [31:0] Q63_375;
wire signed [31:0] Q64_94;
wire signed [31:0] Q64_117;
wire signed [31:0] Q64_132;
wire signed [31:0] Q64_192;
wire signed [31:0] Q64_280;
wire signed [31:0] Q64_352;
wire signed [31:0] Q64_376;
wire signed [31:0] Q65_95;
wire signed [31:0] Q65_118;
wire signed [31:0] Q65_133;
wire signed [31:0] Q65_169;
wire signed [31:0] Q65_281;
wire signed [31:0] Q65_353;
wire signed [31:0] Q65_377;
wire signed [31:0] Q66_96;
wire signed [31:0] Q66_119;
wire signed [31:0] Q66_134;
wire signed [31:0] Q66_170;
wire signed [31:0] Q66_282;
wire signed [31:0] Q66_354;
wire signed [31:0] Q66_378;
wire signed [31:0] Q67_73;
wire signed [31:0] Q67_120;
wire signed [31:0] Q67_135;
wire signed [31:0] Q67_171;
wire signed [31:0] Q67_283;
wire signed [31:0] Q67_355;
wire signed [31:0] Q67_379;
wire signed [31:0] Q68_74;
wire signed [31:0] Q68_97;
wire signed [31:0] Q68_136;
wire signed [31:0] Q68_172;
wire signed [31:0] Q68_284;
wire signed [31:0] Q68_356;
wire signed [31:0] Q68_380;
wire signed [31:0] Q69_75;
wire signed [31:0] Q69_98;
wire signed [31:0] Q69_137;
wire signed [31:0] Q69_173;
wire signed [31:0] Q69_285;
wire signed [31:0] Q69_357;
wire signed [31:0] Q69_381;
wire signed [31:0] Q70_76;
wire signed [31:0] Q70_99;
wire signed [31:0] Q70_138;
wire signed [31:0] Q70_174;
wire signed [31:0] Q70_286;
wire signed [31:0] Q70_358;
wire signed [31:0] Q70_382;
wire signed [31:0] Q71_77;
wire signed [31:0] Q71_100;
wire signed [31:0] Q71_139;
wire signed [31:0] Q71_175;
wire signed [31:0] Q71_287;
wire signed [31:0] Q71_359;
wire signed [31:0] Q71_383;
wire signed [31:0] Q72_78;
wire signed [31:0] Q72_101;
wire signed [31:0] Q72_140;
wire signed [31:0] Q72_176;
wire signed [31:0] Q72_288;
wire signed [31:0] Q72_360;
wire signed [31:0] Q72_384;
wire signed [31:0] Q73_16;
wire signed [31:0] Q73_60;
wire signed [31:0] Q73_209;
wire signed [31:0] Q73_223;
wire signed [31:0] Q73_361;
wire signed [31:0] Q73_385;
wire signed [31:0] Q74_17;
wire signed [31:0] Q74_61;
wire signed [31:0] Q74_210;
wire signed [31:0] Q74_224;
wire signed [31:0] Q74_362;
wire signed [31:0] Q74_386;
wire signed [31:0] Q75_18;
wire signed [31:0] Q75_62;
wire signed [31:0] Q75_211;
wire signed [31:0] Q75_225;
wire signed [31:0] Q75_363;
wire signed [31:0] Q75_387;
wire signed [31:0] Q76_19;
wire signed [31:0] Q76_63;
wire signed [31:0] Q76_212;
wire signed [31:0] Q76_226;
wire signed [31:0] Q76_364;
wire signed [31:0] Q76_388;
wire signed [31:0] Q77_20;
wire signed [31:0] Q77_64;
wire signed [31:0] Q77_213;
wire signed [31:0] Q77_227;
wire signed [31:0] Q77_365;
wire signed [31:0] Q77_389;
wire signed [31:0] Q78_21;
wire signed [31:0] Q78_65;
wire signed [31:0] Q78_214;
wire signed [31:0] Q78_228;
wire signed [31:0] Q78_366;
wire signed [31:0] Q78_390;
wire signed [31:0] Q79_22;
wire signed [31:0] Q79_66;
wire signed [31:0] Q79_215;
wire signed [31:0] Q79_229;
wire signed [31:0] Q79_367;
wire signed [31:0] Q79_391;
wire signed [31:0] Q80_23;
wire signed [31:0] Q80_67;
wire signed [31:0] Q80_216;
wire signed [31:0] Q80_230;
wire signed [31:0] Q80_368;
wire signed [31:0] Q80_392;
wire signed [31:0] Q81_24;
wire signed [31:0] Q81_68;
wire signed [31:0] Q81_193;
wire signed [31:0] Q81_231;
wire signed [31:0] Q81_369;
wire signed [31:0] Q81_393;
wire signed [31:0] Q82_1;
wire signed [31:0] Q82_69;
wire signed [31:0] Q82_194;
wire signed [31:0] Q82_232;
wire signed [31:0] Q82_370;
wire signed [31:0] Q82_394;
wire signed [31:0] Q83_2;
wire signed [31:0] Q83_70;
wire signed [31:0] Q83_195;
wire signed [31:0] Q83_233;
wire signed [31:0] Q83_371;
wire signed [31:0] Q83_395;
wire signed [31:0] Q84_3;
wire signed [31:0] Q84_71;
wire signed [31:0] Q84_196;
wire signed [31:0] Q84_234;
wire signed [31:0] Q84_372;
wire signed [31:0] Q84_396;
wire signed [31:0] Q85_4;
wire signed [31:0] Q85_72;
wire signed [31:0] Q85_197;
wire signed [31:0] Q85_235;
wire signed [31:0] Q85_373;
wire signed [31:0] Q85_397;
wire signed [31:0] Q86_5;
wire signed [31:0] Q86_49;
wire signed [31:0] Q86_198;
wire signed [31:0] Q86_236;
wire signed [31:0] Q86_374;
wire signed [31:0] Q86_398;
wire signed [31:0] Q87_6;
wire signed [31:0] Q87_50;
wire signed [31:0] Q87_199;
wire signed [31:0] Q87_237;
wire signed [31:0] Q87_375;
wire signed [31:0] Q87_399;
wire signed [31:0] Q88_7;
wire signed [31:0] Q88_51;
wire signed [31:0] Q88_200;
wire signed [31:0] Q88_238;
wire signed [31:0] Q88_376;
wire signed [31:0] Q88_400;
wire signed [31:0] Q89_8;
wire signed [31:0] Q89_52;
wire signed [31:0] Q89_201;
wire signed [31:0] Q89_239;
wire signed [31:0] Q89_377;
wire signed [31:0] Q89_401;
wire signed [31:0] Q90_9;
wire signed [31:0] Q90_53;
wire signed [31:0] Q90_202;
wire signed [31:0] Q90_240;
wire signed [31:0] Q90_378;
wire signed [31:0] Q90_402;
wire signed [31:0] Q91_10;
wire signed [31:0] Q91_54;
wire signed [31:0] Q91_203;
wire signed [31:0] Q91_217;
wire signed [31:0] Q91_379;
wire signed [31:0] Q91_403;
wire signed [31:0] Q92_11;
wire signed [31:0] Q92_55;
wire signed [31:0] Q92_204;
wire signed [31:0] Q92_218;
wire signed [31:0] Q92_380;
wire signed [31:0] Q92_404;
wire signed [31:0] Q93_12;
wire signed [31:0] Q93_56;
wire signed [31:0] Q93_205;
wire signed [31:0] Q93_219;
wire signed [31:0] Q93_381;
wire signed [31:0] Q93_405;
wire signed [31:0] Q94_13;
wire signed [31:0] Q94_57;
wire signed [31:0] Q94_206;
wire signed [31:0] Q94_220;
wire signed [31:0] Q94_382;
wire signed [31:0] Q94_406;
wire signed [31:0] Q95_14;
wire signed [31:0] Q95_58;
wire signed [31:0] Q95_207;
wire signed [31:0] Q95_221;
wire signed [31:0] Q95_383;
wire signed [31:0] Q95_407;
wire signed [31:0] Q96_15;
wire signed [31:0] Q96_59;
wire signed [31:0] Q96_208;
wire signed [31:0] Q96_222;
wire signed [31:0] Q96_384;
wire signed [31:0] Q96_408;
wire signed [31:0] Q97_58;
wire signed [31:0] Q97_166;
wire signed [31:0] Q97_227;
wire signed [31:0] Q97_259;
wire signed [31:0] Q97_385;
wire signed [31:0] Q97_409;
wire signed [31:0] Q98_59;
wire signed [31:0] Q98_167;
wire signed [31:0] Q98_228;
wire signed [31:0] Q98_260;
wire signed [31:0] Q98_386;
wire signed [31:0] Q98_410;
wire signed [31:0] Q99_60;
wire signed [31:0] Q99_168;
wire signed [31:0] Q99_229;
wire signed [31:0] Q99_261;
wire signed [31:0] Q99_387;
wire signed [31:0] Q99_411;
wire signed [31:0] Q100_61;
wire signed [31:0] Q100_145;
wire signed [31:0] Q100_230;
wire signed [31:0] Q100_262;
wire signed [31:0] Q100_388;
wire signed [31:0] Q100_412;
wire signed [31:0] Q101_62;
wire signed [31:0] Q101_146;
wire signed [31:0] Q101_231;
wire signed [31:0] Q101_263;
wire signed [31:0] Q101_389;
wire signed [31:0] Q101_413;
wire signed [31:0] Q102_63;
wire signed [31:0] Q102_147;
wire signed [31:0] Q102_232;
wire signed [31:0] Q102_264;
wire signed [31:0] Q102_390;
wire signed [31:0] Q102_414;
wire signed [31:0] Q103_64;
wire signed [31:0] Q103_148;
wire signed [31:0] Q103_233;
wire signed [31:0] Q103_241;
wire signed [31:0] Q103_391;
wire signed [31:0] Q103_415;
wire signed [31:0] Q104_65;
wire signed [31:0] Q104_149;
wire signed [31:0] Q104_234;
wire signed [31:0] Q104_242;
wire signed [31:0] Q104_392;
wire signed [31:0] Q104_416;
wire signed [31:0] Q105_66;
wire signed [31:0] Q105_150;
wire signed [31:0] Q105_235;
wire signed [31:0] Q105_243;
wire signed [31:0] Q105_393;
wire signed [31:0] Q105_417;
wire signed [31:0] Q106_67;
wire signed [31:0] Q106_151;
wire signed [31:0] Q106_236;
wire signed [31:0] Q106_244;
wire signed [31:0] Q106_394;
wire signed [31:0] Q106_418;
wire signed [31:0] Q107_68;
wire signed [31:0] Q107_152;
wire signed [31:0] Q107_237;
wire signed [31:0] Q107_245;
wire signed [31:0] Q107_395;
wire signed [31:0] Q107_419;
wire signed [31:0] Q108_69;
wire signed [31:0] Q108_153;
wire signed [31:0] Q108_238;
wire signed [31:0] Q108_246;
wire signed [31:0] Q108_396;
wire signed [31:0] Q108_420;
wire signed [31:0] Q109_70;
wire signed [31:0] Q109_154;
wire signed [31:0] Q109_239;
wire signed [31:0] Q109_247;
wire signed [31:0] Q109_397;
wire signed [31:0] Q109_421;
wire signed [31:0] Q110_71;
wire signed [31:0] Q110_155;
wire signed [31:0] Q110_240;
wire signed [31:0] Q110_248;
wire signed [31:0] Q110_398;
wire signed [31:0] Q110_422;
wire signed [31:0] Q111_72;
wire signed [31:0] Q111_156;
wire signed [31:0] Q111_217;
wire signed [31:0] Q111_249;
wire signed [31:0] Q111_399;
wire signed [31:0] Q111_423;
wire signed [31:0] Q112_49;
wire signed [31:0] Q112_157;
wire signed [31:0] Q112_218;
wire signed [31:0] Q112_250;
wire signed [31:0] Q112_400;
wire signed [31:0] Q112_424;
wire signed [31:0] Q113_50;
wire signed [31:0] Q113_158;
wire signed [31:0] Q113_219;
wire signed [31:0] Q113_251;
wire signed [31:0] Q113_401;
wire signed [31:0] Q113_425;
wire signed [31:0] Q114_51;
wire signed [31:0] Q114_159;
wire signed [31:0] Q114_220;
wire signed [31:0] Q114_252;
wire signed [31:0] Q114_402;
wire signed [31:0] Q114_426;
wire signed [31:0] Q115_52;
wire signed [31:0] Q115_160;
wire signed [31:0] Q115_221;
wire signed [31:0] Q115_253;
wire signed [31:0] Q115_403;
wire signed [31:0] Q115_427;
wire signed [31:0] Q116_53;
wire signed [31:0] Q116_161;
wire signed [31:0] Q116_222;
wire signed [31:0] Q116_254;
wire signed [31:0] Q116_404;
wire signed [31:0] Q116_428;
wire signed [31:0] Q117_54;
wire signed [31:0] Q117_162;
wire signed [31:0] Q117_223;
wire signed [31:0] Q117_255;
wire signed [31:0] Q117_405;
wire signed [31:0] Q117_429;
wire signed [31:0] Q118_55;
wire signed [31:0] Q118_163;
wire signed [31:0] Q118_224;
wire signed [31:0] Q118_256;
wire signed [31:0] Q118_406;
wire signed [31:0] Q118_430;
wire signed [31:0] Q119_56;
wire signed [31:0] Q119_164;
wire signed [31:0] Q119_225;
wire signed [31:0] Q119_257;
wire signed [31:0] Q119_407;
wire signed [31:0] Q119_431;
wire signed [31:0] Q120_57;
wire signed [31:0] Q120_165;
wire signed [31:0] Q120_226;
wire signed [31:0] Q120_258;
wire signed [31:0] Q120_408;
wire signed [31:0] Q120_432;
wire signed [31:0] Q121_108;
wire signed [31:0] Q121_131;
wire signed [31:0] Q121_189;
wire signed [31:0] Q121_284;
wire signed [31:0] Q121_289;
wire signed [31:0] Q121_409;
wire signed [31:0] Q121_433;
wire signed [31:0] Q122_109;
wire signed [31:0] Q122_132;
wire signed [31:0] Q122_190;
wire signed [31:0] Q122_285;
wire signed [31:0] Q122_290;
wire signed [31:0] Q122_410;
wire signed [31:0] Q122_434;
wire signed [31:0] Q123_110;
wire signed [31:0] Q123_133;
wire signed [31:0] Q123_191;
wire signed [31:0] Q123_286;
wire signed [31:0] Q123_291;
wire signed [31:0] Q123_411;
wire signed [31:0] Q123_435;
wire signed [31:0] Q124_111;
wire signed [31:0] Q124_134;
wire signed [31:0] Q124_192;
wire signed [31:0] Q124_287;
wire signed [31:0] Q124_292;
wire signed [31:0] Q124_412;
wire signed [31:0] Q124_436;
wire signed [31:0] Q125_112;
wire signed [31:0] Q125_135;
wire signed [31:0] Q125_169;
wire signed [31:0] Q125_288;
wire signed [31:0] Q125_293;
wire signed [31:0] Q125_413;
wire signed [31:0] Q125_437;
wire signed [31:0] Q126_113;
wire signed [31:0] Q126_136;
wire signed [31:0] Q126_170;
wire signed [31:0] Q126_265;
wire signed [31:0] Q126_294;
wire signed [31:0] Q126_414;
wire signed [31:0] Q126_438;
wire signed [31:0] Q127_114;
wire signed [31:0] Q127_137;
wire signed [31:0] Q127_171;
wire signed [31:0] Q127_266;
wire signed [31:0] Q127_295;
wire signed [31:0] Q127_415;
wire signed [31:0] Q127_439;
wire signed [31:0] Q128_115;
wire signed [31:0] Q128_138;
wire signed [31:0] Q128_172;
wire signed [31:0] Q128_267;
wire signed [31:0] Q128_296;
wire signed [31:0] Q128_416;
wire signed [31:0] Q128_440;
wire signed [31:0] Q129_116;
wire signed [31:0] Q129_139;
wire signed [31:0] Q129_173;
wire signed [31:0] Q129_268;
wire signed [31:0] Q129_297;
wire signed [31:0] Q129_417;
wire signed [31:0] Q129_441;
wire signed [31:0] Q130_117;
wire signed [31:0] Q130_140;
wire signed [31:0] Q130_174;
wire signed [31:0] Q130_269;
wire signed [31:0] Q130_298;
wire signed [31:0] Q130_418;
wire signed [31:0] Q130_442;
wire signed [31:0] Q131_118;
wire signed [31:0] Q131_141;
wire signed [31:0] Q131_175;
wire signed [31:0] Q131_270;
wire signed [31:0] Q131_299;
wire signed [31:0] Q131_419;
wire signed [31:0] Q131_443;
wire signed [31:0] Q132_119;
wire signed [31:0] Q132_142;
wire signed [31:0] Q132_176;
wire signed [31:0] Q132_271;
wire signed [31:0] Q132_300;
wire signed [31:0] Q132_420;
wire signed [31:0] Q132_444;
wire signed [31:0] Q133_120;
wire signed [31:0] Q133_143;
wire signed [31:0] Q133_177;
wire signed [31:0] Q133_272;
wire signed [31:0] Q133_301;
wire signed [31:0] Q133_421;
wire signed [31:0] Q133_445;
wire signed [31:0] Q134_97;
wire signed [31:0] Q134_144;
wire signed [31:0] Q134_178;
wire signed [31:0] Q134_273;
wire signed [31:0] Q134_302;
wire signed [31:0] Q134_422;
wire signed [31:0] Q134_446;
wire signed [31:0] Q135_98;
wire signed [31:0] Q135_121;
wire signed [31:0] Q135_179;
wire signed [31:0] Q135_274;
wire signed [31:0] Q135_303;
wire signed [31:0] Q135_423;
wire signed [31:0] Q135_447;
wire signed [31:0] Q136_99;
wire signed [31:0] Q136_122;
wire signed [31:0] Q136_180;
wire signed [31:0] Q136_275;
wire signed [31:0] Q136_304;
wire signed [31:0] Q136_424;
wire signed [31:0] Q136_448;
wire signed [31:0] Q137_100;
wire signed [31:0] Q137_123;
wire signed [31:0] Q137_181;
wire signed [31:0] Q137_276;
wire signed [31:0] Q137_305;
wire signed [31:0] Q137_425;
wire signed [31:0] Q137_449;
wire signed [31:0] Q138_101;
wire signed [31:0] Q138_124;
wire signed [31:0] Q138_182;
wire signed [31:0] Q138_277;
wire signed [31:0] Q138_306;
wire signed [31:0] Q138_426;
wire signed [31:0] Q138_450;
wire signed [31:0] Q139_102;
wire signed [31:0] Q139_125;
wire signed [31:0] Q139_183;
wire signed [31:0] Q139_278;
wire signed [31:0] Q139_307;
wire signed [31:0] Q139_427;
wire signed [31:0] Q139_451;
wire signed [31:0] Q140_103;
wire signed [31:0] Q140_126;
wire signed [31:0] Q140_184;
wire signed [31:0] Q140_279;
wire signed [31:0] Q140_308;
wire signed [31:0] Q140_428;
wire signed [31:0] Q140_452;
wire signed [31:0] Q141_104;
wire signed [31:0] Q141_127;
wire signed [31:0] Q141_185;
wire signed [31:0] Q141_280;
wire signed [31:0] Q141_309;
wire signed [31:0] Q141_429;
wire signed [31:0] Q141_453;
wire signed [31:0] Q142_105;
wire signed [31:0] Q142_128;
wire signed [31:0] Q142_186;
wire signed [31:0] Q142_281;
wire signed [31:0] Q142_310;
wire signed [31:0] Q142_430;
wire signed [31:0] Q142_454;
wire signed [31:0] Q143_106;
wire signed [31:0] Q143_129;
wire signed [31:0] Q143_187;
wire signed [31:0] Q143_282;
wire signed [31:0] Q143_311;
wire signed [31:0] Q143_431;
wire signed [31:0] Q143_455;
wire signed [31:0] Q144_107;
wire signed [31:0] Q144_130;
wire signed [31:0] Q144_188;
wire signed [31:0] Q144_283;
wire signed [31:0] Q144_312;
wire signed [31:0] Q144_432;
wire signed [31:0] Q144_456;
wire signed [31:0] Q145_72;
wire signed [31:0] Q145_86;
wire signed [31:0] Q145_220;
wire signed [31:0] Q145_245;
wire signed [31:0] Q145_433;
wire signed [31:0] Q145_457;
wire signed [31:0] Q146_49;
wire signed [31:0] Q146_87;
wire signed [31:0] Q146_221;
wire signed [31:0] Q146_246;
wire signed [31:0] Q146_434;
wire signed [31:0] Q146_458;
wire signed [31:0] Q147_50;
wire signed [31:0] Q147_88;
wire signed [31:0] Q147_222;
wire signed [31:0] Q147_247;
wire signed [31:0] Q147_435;
wire signed [31:0] Q147_459;
wire signed [31:0] Q148_51;
wire signed [31:0] Q148_89;
wire signed [31:0] Q148_223;
wire signed [31:0] Q148_248;
wire signed [31:0] Q148_436;
wire signed [31:0] Q148_460;
wire signed [31:0] Q149_52;
wire signed [31:0] Q149_90;
wire signed [31:0] Q149_224;
wire signed [31:0] Q149_249;
wire signed [31:0] Q149_437;
wire signed [31:0] Q149_461;
wire signed [31:0] Q150_53;
wire signed [31:0] Q150_91;
wire signed [31:0] Q150_225;
wire signed [31:0] Q150_250;
wire signed [31:0] Q150_438;
wire signed [31:0] Q150_462;
wire signed [31:0] Q151_54;
wire signed [31:0] Q151_92;
wire signed [31:0] Q151_226;
wire signed [31:0] Q151_251;
wire signed [31:0] Q151_439;
wire signed [31:0] Q151_463;
wire signed [31:0] Q152_55;
wire signed [31:0] Q152_93;
wire signed [31:0] Q152_227;
wire signed [31:0] Q152_252;
wire signed [31:0] Q152_440;
wire signed [31:0] Q152_464;
wire signed [31:0] Q153_56;
wire signed [31:0] Q153_94;
wire signed [31:0] Q153_228;
wire signed [31:0] Q153_253;
wire signed [31:0] Q153_441;
wire signed [31:0] Q153_465;
wire signed [31:0] Q154_57;
wire signed [31:0] Q154_95;
wire signed [31:0] Q154_229;
wire signed [31:0] Q154_254;
wire signed [31:0] Q154_442;
wire signed [31:0] Q154_466;
wire signed [31:0] Q155_58;
wire signed [31:0] Q155_96;
wire signed [31:0] Q155_230;
wire signed [31:0] Q155_255;
wire signed [31:0] Q155_443;
wire signed [31:0] Q155_467;
wire signed [31:0] Q156_59;
wire signed [31:0] Q156_73;
wire signed [31:0] Q156_231;
wire signed [31:0] Q156_256;
wire signed [31:0] Q156_444;
wire signed [31:0] Q156_468;
wire signed [31:0] Q157_60;
wire signed [31:0] Q157_74;
wire signed [31:0] Q157_232;
wire signed [31:0] Q157_257;
wire signed [31:0] Q157_445;
wire signed [31:0] Q157_469;
wire signed [31:0] Q158_61;
wire signed [31:0] Q158_75;
wire signed [31:0] Q158_233;
wire signed [31:0] Q158_258;
wire signed [31:0] Q158_446;
wire signed [31:0] Q158_470;
wire signed [31:0] Q159_62;
wire signed [31:0] Q159_76;
wire signed [31:0] Q159_234;
wire signed [31:0] Q159_259;
wire signed [31:0] Q159_447;
wire signed [31:0] Q159_471;
wire signed [31:0] Q160_63;
wire signed [31:0] Q160_77;
wire signed [31:0] Q160_235;
wire signed [31:0] Q160_260;
wire signed [31:0] Q160_448;
wire signed [31:0] Q160_472;
wire signed [31:0] Q161_64;
wire signed [31:0] Q161_78;
wire signed [31:0] Q161_236;
wire signed [31:0] Q161_261;
wire signed [31:0] Q161_449;
wire signed [31:0] Q161_473;
wire signed [31:0] Q162_65;
wire signed [31:0] Q162_79;
wire signed [31:0] Q162_237;
wire signed [31:0] Q162_262;
wire signed [31:0] Q162_450;
wire signed [31:0] Q162_474;
wire signed [31:0] Q163_66;
wire signed [31:0] Q163_80;
wire signed [31:0] Q163_238;
wire signed [31:0] Q163_263;
wire signed [31:0] Q163_451;
wire signed [31:0] Q163_475;
wire signed [31:0] Q164_67;
wire signed [31:0] Q164_81;
wire signed [31:0] Q164_239;
wire signed [31:0] Q164_264;
wire signed [31:0] Q164_452;
wire signed [31:0] Q164_476;
wire signed [31:0] Q165_68;
wire signed [31:0] Q165_82;
wire signed [31:0] Q165_240;
wire signed [31:0] Q165_241;
wire signed [31:0] Q165_453;
wire signed [31:0] Q165_477;
wire signed [31:0] Q166_69;
wire signed [31:0] Q166_83;
wire signed [31:0] Q166_217;
wire signed [31:0] Q166_242;
wire signed [31:0] Q166_454;
wire signed [31:0] Q166_478;
wire signed [31:0] Q167_70;
wire signed [31:0] Q167_84;
wire signed [31:0] Q167_218;
wire signed [31:0] Q167_243;
wire signed [31:0] Q167_455;
wire signed [31:0] Q167_479;
wire signed [31:0] Q168_71;
wire signed [31:0] Q168_85;
wire signed [31:0] Q168_219;
wire signed [31:0] Q168_244;
wire signed [31:0] Q168_456;
wire signed [31:0] Q168_480;
wire signed [31:0] Q169_27;
wire signed [31:0] Q169_67;
wire signed [31:0] Q169_145;
wire signed [31:0] Q169_228;
wire signed [31:0] Q169_457;
wire signed [31:0] Q169_481;
wire signed [31:0] Q170_28;
wire signed [31:0] Q170_68;
wire signed [31:0] Q170_146;
wire signed [31:0] Q170_229;
wire signed [31:0] Q170_458;
wire signed [31:0] Q170_482;
wire signed [31:0] Q171_29;
wire signed [31:0] Q171_69;
wire signed [31:0] Q171_147;
wire signed [31:0] Q171_230;
wire signed [31:0] Q171_459;
wire signed [31:0] Q171_483;
wire signed [31:0] Q172_30;
wire signed [31:0] Q172_70;
wire signed [31:0] Q172_148;
wire signed [31:0] Q172_231;
wire signed [31:0] Q172_460;
wire signed [31:0] Q172_484;
wire signed [31:0] Q173_31;
wire signed [31:0] Q173_71;
wire signed [31:0] Q173_149;
wire signed [31:0] Q173_232;
wire signed [31:0] Q173_461;
wire signed [31:0] Q173_485;
wire signed [31:0] Q174_32;
wire signed [31:0] Q174_72;
wire signed [31:0] Q174_150;
wire signed [31:0] Q174_233;
wire signed [31:0] Q174_462;
wire signed [31:0] Q174_486;
wire signed [31:0] Q175_33;
wire signed [31:0] Q175_49;
wire signed [31:0] Q175_151;
wire signed [31:0] Q175_234;
wire signed [31:0] Q175_463;
wire signed [31:0] Q175_487;
wire signed [31:0] Q176_34;
wire signed [31:0] Q176_50;
wire signed [31:0] Q176_152;
wire signed [31:0] Q176_235;
wire signed [31:0] Q176_464;
wire signed [31:0] Q176_488;
wire signed [31:0] Q177_35;
wire signed [31:0] Q177_51;
wire signed [31:0] Q177_153;
wire signed [31:0] Q177_236;
wire signed [31:0] Q177_465;
wire signed [31:0] Q177_489;
wire signed [31:0] Q178_36;
wire signed [31:0] Q178_52;
wire signed [31:0] Q178_154;
wire signed [31:0] Q178_237;
wire signed [31:0] Q178_466;
wire signed [31:0] Q178_490;
wire signed [31:0] Q179_37;
wire signed [31:0] Q179_53;
wire signed [31:0] Q179_155;
wire signed [31:0] Q179_238;
wire signed [31:0] Q179_467;
wire signed [31:0] Q179_491;
wire signed [31:0] Q180_38;
wire signed [31:0] Q180_54;
wire signed [31:0] Q180_156;
wire signed [31:0] Q180_239;
wire signed [31:0] Q180_468;
wire signed [31:0] Q180_492;
wire signed [31:0] Q181_39;
wire signed [31:0] Q181_55;
wire signed [31:0] Q181_157;
wire signed [31:0] Q181_240;
wire signed [31:0] Q181_469;
wire signed [31:0] Q181_493;
wire signed [31:0] Q182_40;
wire signed [31:0] Q182_56;
wire signed [31:0] Q182_158;
wire signed [31:0] Q182_217;
wire signed [31:0] Q182_470;
wire signed [31:0] Q182_494;
wire signed [31:0] Q183_41;
wire signed [31:0] Q183_57;
wire signed [31:0] Q183_159;
wire signed [31:0] Q183_218;
wire signed [31:0] Q183_471;
wire signed [31:0] Q183_495;
wire signed [31:0] Q184_42;
wire signed [31:0] Q184_58;
wire signed [31:0] Q184_160;
wire signed [31:0] Q184_219;
wire signed [31:0] Q184_472;
wire signed [31:0] Q184_496;
wire signed [31:0] Q185_43;
wire signed [31:0] Q185_59;
wire signed [31:0] Q185_161;
wire signed [31:0] Q185_220;
wire signed [31:0] Q185_473;
wire signed [31:0] Q185_497;
wire signed [31:0] Q186_44;
wire signed [31:0] Q186_60;
wire signed [31:0] Q186_162;
wire signed [31:0] Q186_221;
wire signed [31:0] Q186_474;
wire signed [31:0] Q186_498;
wire signed [31:0] Q187_45;
wire signed [31:0] Q187_61;
wire signed [31:0] Q187_163;
wire signed [31:0] Q187_222;
wire signed [31:0] Q187_475;
wire signed [31:0] Q187_499;
wire signed [31:0] Q188_46;
wire signed [31:0] Q188_62;
wire signed [31:0] Q188_164;
wire signed [31:0] Q188_223;
wire signed [31:0] Q188_476;
wire signed [31:0] Q188_500;
wire signed [31:0] Q189_47;
wire signed [31:0] Q189_63;
wire signed [31:0] Q189_165;
wire signed [31:0] Q189_224;
wire signed [31:0] Q189_477;
wire signed [31:0] Q189_501;
wire signed [31:0] Q190_48;
wire signed [31:0] Q190_64;
wire signed [31:0] Q190_166;
wire signed [31:0] Q190_225;
wire signed [31:0] Q190_478;
wire signed [31:0] Q190_502;
wire signed [31:0] Q191_25;
wire signed [31:0] Q191_65;
wire signed [31:0] Q191_167;
wire signed [31:0] Q191_226;
wire signed [31:0] Q191_479;
wire signed [31:0] Q191_503;
wire signed [31:0] Q192_26;
wire signed [31:0] Q192_66;
wire signed [31:0] Q192_168;
wire signed [31:0] Q192_227;
wire signed [31:0] Q192_480;
wire signed [31:0] Q192_504;
wire signed [31:0] Q193_4;
wire signed [31:0] Q193_117;
wire signed [31:0] Q193_127;
wire signed [31:0] Q193_179;
wire signed [31:0] Q193_277;
wire signed [31:0] Q193_481;
wire signed [31:0] Q193_505;
wire signed [31:0] Q194_5;
wire signed [31:0] Q194_118;
wire signed [31:0] Q194_128;
wire signed [31:0] Q194_180;
wire signed [31:0] Q194_278;
wire signed [31:0] Q194_482;
wire signed [31:0] Q194_506;
wire signed [31:0] Q195_6;
wire signed [31:0] Q195_119;
wire signed [31:0] Q195_129;
wire signed [31:0] Q195_181;
wire signed [31:0] Q195_279;
wire signed [31:0] Q195_483;
wire signed [31:0] Q195_507;
wire signed [31:0] Q196_7;
wire signed [31:0] Q196_120;
wire signed [31:0] Q196_130;
wire signed [31:0] Q196_182;
wire signed [31:0] Q196_280;
wire signed [31:0] Q196_484;
wire signed [31:0] Q196_508;
wire signed [31:0] Q197_8;
wire signed [31:0] Q197_97;
wire signed [31:0] Q197_131;
wire signed [31:0] Q197_183;
wire signed [31:0] Q197_281;
wire signed [31:0] Q197_485;
wire signed [31:0] Q197_509;
wire signed [31:0] Q198_9;
wire signed [31:0] Q198_98;
wire signed [31:0] Q198_132;
wire signed [31:0] Q198_184;
wire signed [31:0] Q198_282;
wire signed [31:0] Q198_486;
wire signed [31:0] Q198_510;
wire signed [31:0] Q199_10;
wire signed [31:0] Q199_99;
wire signed [31:0] Q199_133;
wire signed [31:0] Q199_185;
wire signed [31:0] Q199_283;
wire signed [31:0] Q199_487;
wire signed [31:0] Q199_511;
wire signed [31:0] Q200_11;
wire signed [31:0] Q200_100;
wire signed [31:0] Q200_134;
wire signed [31:0] Q200_186;
wire signed [31:0] Q200_284;
wire signed [31:0] Q200_488;
wire signed [31:0] Q200_512;
wire signed [31:0] Q201_12;
wire signed [31:0] Q201_101;
wire signed [31:0] Q201_135;
wire signed [31:0] Q201_187;
wire signed [31:0] Q201_285;
wire signed [31:0] Q201_489;
wire signed [31:0] Q201_513;
wire signed [31:0] Q202_13;
wire signed [31:0] Q202_102;
wire signed [31:0] Q202_136;
wire signed [31:0] Q202_188;
wire signed [31:0] Q202_286;
wire signed [31:0] Q202_490;
wire signed [31:0] Q202_514;
wire signed [31:0] Q203_14;
wire signed [31:0] Q203_103;
wire signed [31:0] Q203_137;
wire signed [31:0] Q203_189;
wire signed [31:0] Q203_287;
wire signed [31:0] Q203_491;
wire signed [31:0] Q203_515;
wire signed [31:0] Q204_15;
wire signed [31:0] Q204_104;
wire signed [31:0] Q204_138;
wire signed [31:0] Q204_190;
wire signed [31:0] Q204_288;
wire signed [31:0] Q204_492;
wire signed [31:0] Q204_516;
wire signed [31:0] Q205_16;
wire signed [31:0] Q205_105;
wire signed [31:0] Q205_139;
wire signed [31:0] Q205_191;
wire signed [31:0] Q205_265;
wire signed [31:0] Q205_493;
wire signed [31:0] Q205_517;
wire signed [31:0] Q206_17;
wire signed [31:0] Q206_106;
wire signed [31:0] Q206_140;
wire signed [31:0] Q206_192;
wire signed [31:0] Q206_266;
wire signed [31:0] Q206_494;
wire signed [31:0] Q206_518;
wire signed [31:0] Q207_18;
wire signed [31:0] Q207_107;
wire signed [31:0] Q207_141;
wire signed [31:0] Q207_169;
wire signed [31:0] Q207_267;
wire signed [31:0] Q207_495;
wire signed [31:0] Q207_519;
wire signed [31:0] Q208_19;
wire signed [31:0] Q208_108;
wire signed [31:0] Q208_142;
wire signed [31:0] Q208_170;
wire signed [31:0] Q208_268;
wire signed [31:0] Q208_496;
wire signed [31:0] Q208_520;
wire signed [31:0] Q209_20;
wire signed [31:0] Q209_109;
wire signed [31:0] Q209_143;
wire signed [31:0] Q209_171;
wire signed [31:0] Q209_269;
wire signed [31:0] Q209_497;
wire signed [31:0] Q209_521;
wire signed [31:0] Q210_21;
wire signed [31:0] Q210_110;
wire signed [31:0] Q210_144;
wire signed [31:0] Q210_172;
wire signed [31:0] Q210_270;
wire signed [31:0] Q210_498;
wire signed [31:0] Q210_522;
wire signed [31:0] Q211_22;
wire signed [31:0] Q211_111;
wire signed [31:0] Q211_121;
wire signed [31:0] Q211_173;
wire signed [31:0] Q211_271;
wire signed [31:0] Q211_499;
wire signed [31:0] Q211_523;
wire signed [31:0] Q212_23;
wire signed [31:0] Q212_112;
wire signed [31:0] Q212_122;
wire signed [31:0] Q212_174;
wire signed [31:0] Q212_272;
wire signed [31:0] Q212_500;
wire signed [31:0] Q212_524;
wire signed [31:0] Q213_24;
wire signed [31:0] Q213_113;
wire signed [31:0] Q213_123;
wire signed [31:0] Q213_175;
wire signed [31:0] Q213_273;
wire signed [31:0] Q213_501;
wire signed [31:0] Q213_525;
wire signed [31:0] Q214_1;
wire signed [31:0] Q214_114;
wire signed [31:0] Q214_124;
wire signed [31:0] Q214_176;
wire signed [31:0] Q214_274;
wire signed [31:0] Q214_502;
wire signed [31:0] Q214_526;
wire signed [31:0] Q215_2;
wire signed [31:0] Q215_115;
wire signed [31:0] Q215_125;
wire signed [31:0] Q215_177;
wire signed [31:0] Q215_275;
wire signed [31:0] Q215_503;
wire signed [31:0] Q215_527;
wire signed [31:0] Q216_3;
wire signed [31:0] Q216_116;
wire signed [31:0] Q216_126;
wire signed [31:0] Q216_178;
wire signed [31:0] Q216_276;
wire signed [31:0] Q216_504;
wire signed [31:0] Q216_528;
wire signed [31:0] Q217_144;
wire signed [31:0] Q217_183;
wire signed [31:0] Q217_258;
wire signed [31:0] Q217_283;
wire signed [31:0] Q217_505;
wire signed [31:0] Q217_529;
wire signed [31:0] Q218_121;
wire signed [31:0] Q218_184;
wire signed [31:0] Q218_259;
wire signed [31:0] Q218_284;
wire signed [31:0] Q218_506;
wire signed [31:0] Q218_530;
wire signed [31:0] Q219_122;
wire signed [31:0] Q219_185;
wire signed [31:0] Q219_260;
wire signed [31:0] Q219_285;
wire signed [31:0] Q219_507;
wire signed [31:0] Q219_531;
wire signed [31:0] Q220_123;
wire signed [31:0] Q220_186;
wire signed [31:0] Q220_261;
wire signed [31:0] Q220_286;
wire signed [31:0] Q220_508;
wire signed [31:0] Q220_532;
wire signed [31:0] Q221_124;
wire signed [31:0] Q221_187;
wire signed [31:0] Q221_262;
wire signed [31:0] Q221_287;
wire signed [31:0] Q221_509;
wire signed [31:0] Q221_533;
wire signed [31:0] Q222_125;
wire signed [31:0] Q222_188;
wire signed [31:0] Q222_263;
wire signed [31:0] Q222_288;
wire signed [31:0] Q222_510;
wire signed [31:0] Q222_534;
wire signed [31:0] Q223_126;
wire signed [31:0] Q223_189;
wire signed [31:0] Q223_264;
wire signed [31:0] Q223_265;
wire signed [31:0] Q223_511;
wire signed [31:0] Q223_535;
wire signed [31:0] Q224_127;
wire signed [31:0] Q224_190;
wire signed [31:0] Q224_241;
wire signed [31:0] Q224_266;
wire signed [31:0] Q224_512;
wire signed [31:0] Q224_536;
wire signed [31:0] Q225_128;
wire signed [31:0] Q225_191;
wire signed [31:0] Q225_242;
wire signed [31:0] Q225_267;
wire signed [31:0] Q225_513;
wire signed [31:0] Q225_537;
wire signed [31:0] Q226_129;
wire signed [31:0] Q226_192;
wire signed [31:0] Q226_243;
wire signed [31:0] Q226_268;
wire signed [31:0] Q226_514;
wire signed [31:0] Q226_538;
wire signed [31:0] Q227_130;
wire signed [31:0] Q227_169;
wire signed [31:0] Q227_244;
wire signed [31:0] Q227_269;
wire signed [31:0] Q227_515;
wire signed [31:0] Q227_539;
wire signed [31:0] Q228_131;
wire signed [31:0] Q228_170;
wire signed [31:0] Q228_245;
wire signed [31:0] Q228_270;
wire signed [31:0] Q228_516;
wire signed [31:0] Q228_540;
wire signed [31:0] Q229_132;
wire signed [31:0] Q229_171;
wire signed [31:0] Q229_246;
wire signed [31:0] Q229_271;
wire signed [31:0] Q229_517;
wire signed [31:0] Q229_541;
wire signed [31:0] Q230_133;
wire signed [31:0] Q230_172;
wire signed [31:0] Q230_247;
wire signed [31:0] Q230_272;
wire signed [31:0] Q230_518;
wire signed [31:0] Q230_542;
wire signed [31:0] Q231_134;
wire signed [31:0] Q231_173;
wire signed [31:0] Q231_248;
wire signed [31:0] Q231_273;
wire signed [31:0] Q231_519;
wire signed [31:0] Q231_543;
wire signed [31:0] Q232_135;
wire signed [31:0] Q232_174;
wire signed [31:0] Q232_249;
wire signed [31:0] Q232_274;
wire signed [31:0] Q232_520;
wire signed [31:0] Q232_544;
wire signed [31:0] Q233_136;
wire signed [31:0] Q233_175;
wire signed [31:0] Q233_250;
wire signed [31:0] Q233_275;
wire signed [31:0] Q233_521;
wire signed [31:0] Q233_545;
wire signed [31:0] Q234_137;
wire signed [31:0] Q234_176;
wire signed [31:0] Q234_251;
wire signed [31:0] Q234_276;
wire signed [31:0] Q234_522;
wire signed [31:0] Q234_546;
wire signed [31:0] Q235_138;
wire signed [31:0] Q235_177;
wire signed [31:0] Q235_252;
wire signed [31:0] Q235_277;
wire signed [31:0] Q235_523;
wire signed [31:0] Q235_547;
wire signed [31:0] Q236_139;
wire signed [31:0] Q236_178;
wire signed [31:0] Q236_253;
wire signed [31:0] Q236_278;
wire signed [31:0] Q236_524;
wire signed [31:0] Q236_548;
wire signed [31:0] Q237_140;
wire signed [31:0] Q237_179;
wire signed [31:0] Q237_254;
wire signed [31:0] Q237_279;
wire signed [31:0] Q237_525;
wire signed [31:0] Q237_549;
wire signed [31:0] Q238_141;
wire signed [31:0] Q238_180;
wire signed [31:0] Q238_255;
wire signed [31:0] Q238_280;
wire signed [31:0] Q238_526;
wire signed [31:0] Q238_550;
wire signed [31:0] Q239_142;
wire signed [31:0] Q239_181;
wire signed [31:0] Q239_256;
wire signed [31:0] Q239_281;
wire signed [31:0] Q239_527;
wire signed [31:0] Q239_551;
wire signed [31:0] Q240_143;
wire signed [31:0] Q240_182;
wire signed [31:0] Q240_257;
wire signed [31:0] Q240_282;
wire signed [31:0] Q240_528;
wire signed [31:0] Q240_552;
wire signed [31:0] Q241_50;
wire signed [31:0] Q241_89;
wire signed [31:0] Q241_202;
wire signed [31:0] Q241_229;
wire signed [31:0] Q241_529;
wire signed [31:0] Q241_553;
wire signed [31:0] Q242_51;
wire signed [31:0] Q242_90;
wire signed [31:0] Q242_203;
wire signed [31:0] Q242_230;
wire signed [31:0] Q242_530;
wire signed [31:0] Q242_554;
wire signed [31:0] Q243_52;
wire signed [31:0] Q243_91;
wire signed [31:0] Q243_204;
wire signed [31:0] Q243_231;
wire signed [31:0] Q243_531;
wire signed [31:0] Q243_555;
wire signed [31:0] Q244_53;
wire signed [31:0] Q244_92;
wire signed [31:0] Q244_205;
wire signed [31:0] Q244_232;
wire signed [31:0] Q244_532;
wire signed [31:0] Q244_556;
wire signed [31:0] Q245_54;
wire signed [31:0] Q245_93;
wire signed [31:0] Q245_206;
wire signed [31:0] Q245_233;
wire signed [31:0] Q245_533;
wire signed [31:0] Q245_557;
wire signed [31:0] Q246_55;
wire signed [31:0] Q246_94;
wire signed [31:0] Q246_207;
wire signed [31:0] Q246_234;
wire signed [31:0] Q246_534;
wire signed [31:0] Q246_558;
wire signed [31:0] Q247_56;
wire signed [31:0] Q247_95;
wire signed [31:0] Q247_208;
wire signed [31:0] Q247_235;
wire signed [31:0] Q247_535;
wire signed [31:0] Q247_559;
wire signed [31:0] Q248_57;
wire signed [31:0] Q248_96;
wire signed [31:0] Q248_209;
wire signed [31:0] Q248_236;
wire signed [31:0] Q248_536;
wire signed [31:0] Q248_560;
wire signed [31:0] Q249_58;
wire signed [31:0] Q249_73;
wire signed [31:0] Q249_210;
wire signed [31:0] Q249_237;
wire signed [31:0] Q249_537;
wire signed [31:0] Q249_561;
wire signed [31:0] Q250_59;
wire signed [31:0] Q250_74;
wire signed [31:0] Q250_211;
wire signed [31:0] Q250_238;
wire signed [31:0] Q250_538;
wire signed [31:0] Q250_562;
wire signed [31:0] Q251_60;
wire signed [31:0] Q251_75;
wire signed [31:0] Q251_212;
wire signed [31:0] Q251_239;
wire signed [31:0] Q251_539;
wire signed [31:0] Q251_563;
wire signed [31:0] Q252_61;
wire signed [31:0] Q252_76;
wire signed [31:0] Q252_213;
wire signed [31:0] Q252_240;
wire signed [31:0] Q252_540;
wire signed [31:0] Q252_564;
wire signed [31:0] Q253_62;
wire signed [31:0] Q253_77;
wire signed [31:0] Q253_214;
wire signed [31:0] Q253_217;
wire signed [31:0] Q253_541;
wire signed [31:0] Q253_565;
wire signed [31:0] Q254_63;
wire signed [31:0] Q254_78;
wire signed [31:0] Q254_215;
wire signed [31:0] Q254_218;
wire signed [31:0] Q254_542;
wire signed [31:0] Q254_566;
wire signed [31:0] Q255_64;
wire signed [31:0] Q255_79;
wire signed [31:0] Q255_216;
wire signed [31:0] Q255_219;
wire signed [31:0] Q255_543;
wire signed [31:0] Q255_567;
wire signed [31:0] Q256_65;
wire signed [31:0] Q256_80;
wire signed [31:0] Q256_193;
wire signed [31:0] Q256_220;
wire signed [31:0] Q256_544;
wire signed [31:0] Q256_568;
wire signed [31:0] Q257_66;
wire signed [31:0] Q257_81;
wire signed [31:0] Q257_194;
wire signed [31:0] Q257_221;
wire signed [31:0] Q257_545;
wire signed [31:0] Q257_569;
wire signed [31:0] Q258_67;
wire signed [31:0] Q258_82;
wire signed [31:0] Q258_195;
wire signed [31:0] Q258_222;
wire signed [31:0] Q258_546;
wire signed [31:0] Q258_570;
wire signed [31:0] Q259_68;
wire signed [31:0] Q259_83;
wire signed [31:0] Q259_196;
wire signed [31:0] Q259_223;
wire signed [31:0] Q259_547;
wire signed [31:0] Q259_571;
wire signed [31:0] Q260_69;
wire signed [31:0] Q260_84;
wire signed [31:0] Q260_197;
wire signed [31:0] Q260_224;
wire signed [31:0] Q260_548;
wire signed [31:0] Q260_572;
wire signed [31:0] Q261_70;
wire signed [31:0] Q261_85;
wire signed [31:0] Q261_198;
wire signed [31:0] Q261_225;
wire signed [31:0] Q261_549;
wire signed [31:0] Q261_573;
wire signed [31:0] Q262_71;
wire signed [31:0] Q262_86;
wire signed [31:0] Q262_199;
wire signed [31:0] Q262_226;
wire signed [31:0] Q262_550;
wire signed [31:0] Q262_574;
wire signed [31:0] Q263_72;
wire signed [31:0] Q263_87;
wire signed [31:0] Q263_200;
wire signed [31:0] Q263_227;
wire signed [31:0] Q263_551;
wire signed [31:0] Q263_575;
wire signed [31:0] Q264_49;
wire signed [31:0] Q264_88;
wire signed [31:0] Q264_201;
wire signed [31:0] Q264_228;
wire signed [31:0] Q264_552;
wire signed [31:0] Q264_576;
wire signed [31:0] Q265_11;
wire signed [31:0] Q265_137;
wire signed [31:0] Q265_179;
wire signed [31:0] Q265_271;
wire signed [31:0] Q265_290;
wire signed [31:0] Q265_553;
wire signed [31:0] Q266_12;
wire signed [31:0] Q266_138;
wire signed [31:0] Q266_180;
wire signed [31:0] Q266_272;
wire signed [31:0] Q266_291;
wire signed [31:0] Q266_554;
wire signed [31:0] Q267_13;
wire signed [31:0] Q267_139;
wire signed [31:0] Q267_181;
wire signed [31:0] Q267_273;
wire signed [31:0] Q267_292;
wire signed [31:0] Q267_555;
wire signed [31:0] Q268_14;
wire signed [31:0] Q268_140;
wire signed [31:0] Q268_182;
wire signed [31:0] Q268_274;
wire signed [31:0] Q268_293;
wire signed [31:0] Q268_556;
wire signed [31:0] Q269_15;
wire signed [31:0] Q269_141;
wire signed [31:0] Q269_183;
wire signed [31:0] Q269_275;
wire signed [31:0] Q269_294;
wire signed [31:0] Q269_557;
wire signed [31:0] Q270_16;
wire signed [31:0] Q270_142;
wire signed [31:0] Q270_184;
wire signed [31:0] Q270_276;
wire signed [31:0] Q270_295;
wire signed [31:0] Q270_558;
wire signed [31:0] Q271_17;
wire signed [31:0] Q271_143;
wire signed [31:0] Q271_185;
wire signed [31:0] Q271_277;
wire signed [31:0] Q271_296;
wire signed [31:0] Q271_559;
wire signed [31:0] Q272_18;
wire signed [31:0] Q272_144;
wire signed [31:0] Q272_186;
wire signed [31:0] Q272_278;
wire signed [31:0] Q272_297;
wire signed [31:0] Q272_560;
wire signed [31:0] Q273_19;
wire signed [31:0] Q273_121;
wire signed [31:0] Q273_187;
wire signed [31:0] Q273_279;
wire signed [31:0] Q273_298;
wire signed [31:0] Q273_561;
wire signed [31:0] Q274_20;
wire signed [31:0] Q274_122;
wire signed [31:0] Q274_188;
wire signed [31:0] Q274_280;
wire signed [31:0] Q274_299;
wire signed [31:0] Q274_562;
wire signed [31:0] Q275_21;
wire signed [31:0] Q275_123;
wire signed [31:0] Q275_189;
wire signed [31:0] Q275_281;
wire signed [31:0] Q275_300;
wire signed [31:0] Q275_563;
wire signed [31:0] Q276_22;
wire signed [31:0] Q276_124;
wire signed [31:0] Q276_190;
wire signed [31:0] Q276_282;
wire signed [31:0] Q276_301;
wire signed [31:0] Q276_564;
wire signed [31:0] Q277_23;
wire signed [31:0] Q277_125;
wire signed [31:0] Q277_191;
wire signed [31:0] Q277_283;
wire signed [31:0] Q277_302;
wire signed [31:0] Q277_565;
wire signed [31:0] Q278_24;
wire signed [31:0] Q278_126;
wire signed [31:0] Q278_192;
wire signed [31:0] Q278_284;
wire signed [31:0] Q278_303;
wire signed [31:0] Q278_566;
wire signed [31:0] Q279_1;
wire signed [31:0] Q279_127;
wire signed [31:0] Q279_169;
wire signed [31:0] Q279_285;
wire signed [31:0] Q279_304;
wire signed [31:0] Q279_567;
wire signed [31:0] Q280_2;
wire signed [31:0] Q280_128;
wire signed [31:0] Q280_170;
wire signed [31:0] Q280_286;
wire signed [31:0] Q280_305;
wire signed [31:0] Q280_568;
wire signed [31:0] Q281_3;
wire signed [31:0] Q281_129;
wire signed [31:0] Q281_171;
wire signed [31:0] Q281_287;
wire signed [31:0] Q281_306;
wire signed [31:0] Q281_569;
wire signed [31:0] Q282_4;
wire signed [31:0] Q282_130;
wire signed [31:0] Q282_172;
wire signed [31:0] Q282_288;
wire signed [31:0] Q282_307;
wire signed [31:0] Q282_570;
wire signed [31:0] Q283_5;
wire signed [31:0] Q283_131;
wire signed [31:0] Q283_173;
wire signed [31:0] Q283_265;
wire signed [31:0] Q283_308;
wire signed [31:0] Q283_571;
wire signed [31:0] Q284_6;
wire signed [31:0] Q284_132;
wire signed [31:0] Q284_174;
wire signed [31:0] Q284_266;
wire signed [31:0] Q284_309;
wire signed [31:0] Q284_572;
wire signed [31:0] Q285_7;
wire signed [31:0] Q285_133;
wire signed [31:0] Q285_175;
wire signed [31:0] Q285_267;
wire signed [31:0] Q285_310;
wire signed [31:0] Q285_573;
wire signed [31:0] Q286_8;
wire signed [31:0] Q286_134;
wire signed [31:0] Q286_176;
wire signed [31:0] Q286_268;
wire signed [31:0] Q286_311;
wire signed [31:0] Q286_574;
wire signed [31:0] Q287_9;
wire signed [31:0] Q287_135;
wire signed [31:0] Q287_177;
wire signed [31:0] Q287_269;
wire signed [31:0] Q287_312;
wire signed [31:0] Q287_575;
wire signed [31:0] Q288_10;
wire signed [31:0] Q288_136;
wire signed [31:0] Q288_178;
wire signed [31:0] Q288_270;
wire signed [31:0] Q288_289;
wire signed [31:0] Q288_576;
CNU_6 CNU1(R1_48, R1_67, R1_206, R1_237, R1_290, R1_313, Q1_48, Q1_67, Q1_206, Q1_237, Q1_290, Q1_313, clk );
CNU_6 CNU2(R2_25, R2_68, R2_207, R2_238, R2_291, R2_314, Q2_25, Q2_68, Q2_207, Q2_238, Q2_291, Q2_314, clk );
CNU_6 CNU3(R3_26, R3_69, R3_208, R3_239, R3_292, R3_315, Q3_26, Q3_69, Q3_208, Q3_239, Q3_292, Q3_315, clk );
CNU_6 CNU4(R4_27, R4_70, R4_209, R4_240, R4_293, R4_316, Q4_27, Q4_70, Q4_209, Q4_240, Q4_293, Q4_316, clk );
CNU_6 CNU5(R5_28, R5_71, R5_210, R5_217, R5_294, R5_317, Q5_28, Q5_71, Q5_210, Q5_217, Q5_294, Q5_317, clk );
CNU_6 CNU6(R6_29, R6_72, R6_211, R6_218, R6_295, R6_318, Q6_29, Q6_72, Q6_211, Q6_218, Q6_295, Q6_318, clk );
CNU_6 CNU7(R7_30, R7_49, R7_212, R7_219, R7_296, R7_319, Q7_30, Q7_49, Q7_212, Q7_219, Q7_296, Q7_319, clk );
CNU_6 CNU8(R8_31, R8_50, R8_213, R8_220, R8_297, R8_320, Q8_31, Q8_50, Q8_213, Q8_220, Q8_297, Q8_320, clk );
CNU_6 CNU9(R9_32, R9_51, R9_214, R9_221, R9_298, R9_321, Q9_32, Q9_51, Q9_214, Q9_221, Q9_298, Q9_321, clk );
CNU_6 CNU10(R10_33, R10_52, R10_215, R10_222, R10_299, R10_322, Q10_33, Q10_52, Q10_215, Q10_222, Q10_299, Q10_322, clk );
CNU_6 CNU11(R11_34, R11_53, R11_216, R11_223, R11_300, R11_323, Q11_34, Q11_53, Q11_216, Q11_223, Q11_300, Q11_323, clk );
CNU_6 CNU12(R12_35, R12_54, R12_193, R12_224, R12_301, R12_324, Q12_35, Q12_54, Q12_193, Q12_224, Q12_301, Q12_324, clk );
CNU_6 CNU13(R13_36, R13_55, R13_194, R13_225, R13_302, R13_325, Q13_36, Q13_55, Q13_194, Q13_225, Q13_302, Q13_325, clk );
CNU_6 CNU14(R14_37, R14_56, R14_195, R14_226, R14_303, R14_326, Q14_37, Q14_56, Q14_195, Q14_226, Q14_303, Q14_326, clk );
CNU_6 CNU15(R15_38, R15_57, R15_196, R15_227, R15_304, R15_327, Q15_38, Q15_57, Q15_196, Q15_227, Q15_304, Q15_327, clk );
CNU_6 CNU16(R16_39, R16_58, R16_197, R16_228, R16_305, R16_328, Q16_39, Q16_58, Q16_197, Q16_228, Q16_305, Q16_328, clk );
CNU_6 CNU17(R17_40, R17_59, R17_198, R17_229, R17_306, R17_329, Q17_40, Q17_59, Q17_198, Q17_229, Q17_306, Q17_329, clk );
CNU_6 CNU18(R18_41, R18_60, R18_199, R18_230, R18_307, R18_330, Q18_41, Q18_60, Q18_199, Q18_230, Q18_307, Q18_330, clk );
CNU_6 CNU19(R19_42, R19_61, R19_200, R19_231, R19_308, R19_331, Q19_42, Q19_61, Q19_200, Q19_231, Q19_308, Q19_331, clk );
CNU_6 CNU20(R20_43, R20_62, R20_201, R20_232, R20_309, R20_332, Q20_43, Q20_62, Q20_201, Q20_232, Q20_309, Q20_332, clk );
CNU_6 CNU21(R21_44, R21_63, R21_202, R21_233, R21_310, R21_333, Q21_44, Q21_63, Q21_202, Q21_233, Q21_310, Q21_333, clk );
CNU_6 CNU22(R22_45, R22_64, R22_203, R22_234, R22_311, R22_334, Q22_45, Q22_64, Q22_203, Q22_234, Q22_311, Q22_334, clk );
CNU_6 CNU23(R23_46, R23_65, R23_204, R23_235, R23_312, R23_335, Q23_46, Q23_65, Q23_204, Q23_235, Q23_312, Q23_335, clk );
CNU_6 CNU24(R24_47, R24_66, R24_205, R24_236, R24_289, R24_336, Q24_47, Q24_66, Q24_205, Q24_236, Q24_289, Q24_336, clk );
CNU_7 CNU25(R25_31, R25_126, R25_164, R25_171, R25_268, R25_313, R25_337, Q25_31, Q25_126, Q25_164, Q25_171, Q25_268, Q25_313, Q25_337, clk );
CNU_7 CNU26(R26_32, R26_127, R26_165, R26_172, R26_269, R26_314, R26_338, Q26_32, Q26_127, Q26_165, Q26_172, Q26_269, Q26_314, Q26_338, clk );
CNU_7 CNU27(R27_33, R27_128, R27_166, R27_173, R27_270, R27_315, R27_339, Q27_33, Q27_128, Q27_166, Q27_173, Q27_270, Q27_315, Q27_339, clk );
CNU_7 CNU28(R28_34, R28_129, R28_167, R28_174, R28_271, R28_316, R28_340, Q28_34, Q28_129, Q28_167, Q28_174, Q28_271, Q28_316, Q28_340, clk );
CNU_7 CNU29(R29_35, R29_130, R29_168, R29_175, R29_272, R29_317, R29_341, Q29_35, Q29_130, Q29_168, Q29_175, Q29_272, Q29_317, Q29_341, clk );
CNU_7 CNU30(R30_36, R30_131, R30_145, R30_176, R30_273, R30_318, R30_342, Q30_36, Q30_131, Q30_145, Q30_176, Q30_273, Q30_318, Q30_342, clk );
CNU_7 CNU31(R31_37, R31_132, R31_146, R31_177, R31_274, R31_319, R31_343, Q31_37, Q31_132, Q31_146, Q31_177, Q31_274, Q31_319, Q31_343, clk );
CNU_7 CNU32(R32_38, R32_133, R32_147, R32_178, R32_275, R32_320, R32_344, Q32_38, Q32_133, Q32_147, Q32_178, Q32_275, Q32_320, Q32_344, clk );
CNU_7 CNU33(R33_39, R33_134, R33_148, R33_179, R33_276, R33_321, R33_345, Q33_39, Q33_134, Q33_148, Q33_179, Q33_276, Q33_321, Q33_345, clk );
CNU_7 CNU34(R34_40, R34_135, R34_149, R34_180, R34_277, R34_322, R34_346, Q34_40, Q34_135, Q34_149, Q34_180, Q34_277, Q34_322, Q34_346, clk );
CNU_7 CNU35(R35_41, R35_136, R35_150, R35_181, R35_278, R35_323, R35_347, Q35_41, Q35_136, Q35_150, Q35_181, Q35_278, Q35_323, Q35_347, clk );
CNU_7 CNU36(R36_42, R36_137, R36_151, R36_182, R36_279, R36_324, R36_348, Q36_42, Q36_137, Q36_151, Q36_182, Q36_279, Q36_324, Q36_348, clk );
CNU_7 CNU37(R37_43, R37_138, R37_152, R37_183, R37_280, R37_325, R37_349, Q37_43, Q37_138, Q37_152, Q37_183, Q37_280, Q37_325, Q37_349, clk );
CNU_7 CNU38(R38_44, R38_139, R38_153, R38_184, R38_281, R38_326, R38_350, Q38_44, Q38_139, Q38_153, Q38_184, Q38_281, Q38_326, Q38_350, clk );
CNU_7 CNU39(R39_45, R39_140, R39_154, R39_185, R39_282, R39_327, R39_351, Q39_45, Q39_140, Q39_154, Q39_185, Q39_282, Q39_327, Q39_351, clk );
CNU_7 CNU40(R40_46, R40_141, R40_155, R40_186, R40_283, R40_328, R40_352, Q40_46, Q40_141, Q40_155, Q40_186, Q40_283, Q40_328, Q40_352, clk );
CNU_7 CNU41(R41_47, R41_142, R41_156, R41_187, R41_284, R41_329, R41_353, Q41_47, Q41_142, Q41_156, Q41_187, Q41_284, Q41_329, Q41_353, clk );
CNU_7 CNU42(R42_48, R42_143, R42_157, R42_188, R42_285, R42_330, R42_354, Q42_48, Q42_143, Q42_157, Q42_188, Q42_285, Q42_330, Q42_354, clk );
CNU_7 CNU43(R43_25, R43_144, R43_158, R43_189, R43_286, R43_331, R43_355, Q43_25, Q43_144, Q43_158, Q43_189, Q43_286, Q43_331, Q43_355, clk );
CNU_7 CNU44(R44_26, R44_121, R44_159, R44_190, R44_287, R44_332, R44_356, Q44_26, Q44_121, Q44_159, Q44_190, Q44_287, Q44_332, Q44_356, clk );
CNU_7 CNU45(R45_27, R45_122, R45_160, R45_191, R45_288, R45_333, R45_357, Q45_27, Q45_122, Q45_160, Q45_191, Q45_288, Q45_333, Q45_357, clk );
CNU_7 CNU46(R46_28, R46_123, R46_161, R46_192, R46_265, R46_334, R46_358, Q46_28, Q46_123, Q46_161, Q46_192, Q46_265, Q46_334, Q46_358, clk );
CNU_7 CNU47(R47_29, R47_124, R47_162, R47_169, R47_266, R47_335, R47_359, Q47_29, Q47_124, Q47_162, Q47_169, Q47_266, Q47_335, Q47_359, clk );
CNU_7 CNU48(R48_30, R48_125, R48_163, R48_170, R48_267, R48_336, R48_360, Q48_30, Q48_125, Q48_163, Q48_170, Q48_267, Q48_336, Q48_360, clk );
CNU_7 CNU49(R49_79, R49_102, R49_141, R49_177, R49_265, R49_337, R49_361, Q49_79, Q49_102, Q49_141, Q49_177, Q49_265, Q49_337, Q49_361, clk );
CNU_7 CNU50(R50_80, R50_103, R50_142, R50_178, R50_266, R50_338, R50_362, Q50_80, Q50_103, Q50_142, Q50_178, Q50_266, Q50_338, Q50_362, clk );
CNU_7 CNU51(R51_81, R51_104, R51_143, R51_179, R51_267, R51_339, R51_363, Q51_81, Q51_104, Q51_143, Q51_179, Q51_267, Q51_339, Q51_363, clk );
CNU_7 CNU52(R52_82, R52_105, R52_144, R52_180, R52_268, R52_340, R52_364, Q52_82, Q52_105, Q52_144, Q52_180, Q52_268, Q52_340, Q52_364, clk );
CNU_7 CNU53(R53_83, R53_106, R53_121, R53_181, R53_269, R53_341, R53_365, Q53_83, Q53_106, Q53_121, Q53_181, Q53_269, Q53_341, Q53_365, clk );
CNU_7 CNU54(R54_84, R54_107, R54_122, R54_182, R54_270, R54_342, R54_366, Q54_84, Q54_107, Q54_122, Q54_182, Q54_270, Q54_342, Q54_366, clk );
CNU_7 CNU55(R55_85, R55_108, R55_123, R55_183, R55_271, R55_343, R55_367, Q55_85, Q55_108, Q55_123, Q55_183, Q55_271, Q55_343, Q55_367, clk );
CNU_7 CNU56(R56_86, R56_109, R56_124, R56_184, R56_272, R56_344, R56_368, Q56_86, Q56_109, Q56_124, Q56_184, Q56_272, Q56_344, Q56_368, clk );
CNU_7 CNU57(R57_87, R57_110, R57_125, R57_185, R57_273, R57_345, R57_369, Q57_87, Q57_110, Q57_125, Q57_185, Q57_273, Q57_345, Q57_369, clk );
CNU_7 CNU58(R58_88, R58_111, R58_126, R58_186, R58_274, R58_346, R58_370, Q58_88, Q58_111, Q58_126, Q58_186, Q58_274, Q58_346, Q58_370, clk );
CNU_7 CNU59(R59_89, R59_112, R59_127, R59_187, R59_275, R59_347, R59_371, Q59_89, Q59_112, Q59_127, Q59_187, Q59_275, Q59_347, Q59_371, clk );
CNU_7 CNU60(R60_90, R60_113, R60_128, R60_188, R60_276, R60_348, R60_372, Q60_90, Q60_113, Q60_128, Q60_188, Q60_276, Q60_348, Q60_372, clk );
CNU_7 CNU61(R61_91, R61_114, R61_129, R61_189, R61_277, R61_349, R61_373, Q61_91, Q61_114, Q61_129, Q61_189, Q61_277, Q61_349, Q61_373, clk );
CNU_7 CNU62(R62_92, R62_115, R62_130, R62_190, R62_278, R62_350, R62_374, Q62_92, Q62_115, Q62_130, Q62_190, Q62_278, Q62_350, Q62_374, clk );
CNU_7 CNU63(R63_93, R63_116, R63_131, R63_191, R63_279, R63_351, R63_375, Q63_93, Q63_116, Q63_131, Q63_191, Q63_279, Q63_351, Q63_375, clk );
CNU_7 CNU64(R64_94, R64_117, R64_132, R64_192, R64_280, R64_352, R64_376, Q64_94, Q64_117, Q64_132, Q64_192, Q64_280, Q64_352, Q64_376, clk );
CNU_7 CNU65(R65_95, R65_118, R65_133, R65_169, R65_281, R65_353, R65_377, Q65_95, Q65_118, Q65_133, Q65_169, Q65_281, Q65_353, Q65_377, clk );
CNU_7 CNU66(R66_96, R66_119, R66_134, R66_170, R66_282, R66_354, R66_378, Q66_96, Q66_119, Q66_134, Q66_170, Q66_282, Q66_354, Q66_378, clk );
CNU_7 CNU67(R67_73, R67_120, R67_135, R67_171, R67_283, R67_355, R67_379, Q67_73, Q67_120, Q67_135, Q67_171, Q67_283, Q67_355, Q67_379, clk );
CNU_7 CNU68(R68_74, R68_97, R68_136, R68_172, R68_284, R68_356, R68_380, Q68_74, Q68_97, Q68_136, Q68_172, Q68_284, Q68_356, Q68_380, clk );
CNU_7 CNU69(R69_75, R69_98, R69_137, R69_173, R69_285, R69_357, R69_381, Q69_75, Q69_98, Q69_137, Q69_173, Q69_285, Q69_357, Q69_381, clk );
CNU_7 CNU70(R70_76, R70_99, R70_138, R70_174, R70_286, R70_358, R70_382, Q70_76, Q70_99, Q70_138, Q70_174, Q70_286, Q70_358, Q70_382, clk );
CNU_7 CNU71(R71_77, R71_100, R71_139, R71_175, R71_287, R71_359, R71_383, Q71_77, Q71_100, Q71_139, Q71_175, Q71_287, Q71_359, Q71_383, clk );
CNU_7 CNU72(R72_78, R72_101, R72_140, R72_176, R72_288, R72_360, R72_384, Q72_78, Q72_101, Q72_140, Q72_176, Q72_288, Q72_360, Q72_384, clk );
CNU_6 CNU73(R73_16, R73_60, R73_209, R73_223, R73_361, R73_385, Q73_16, Q73_60, Q73_209, Q73_223, Q73_361, Q73_385, clk );
CNU_6 CNU74(R74_17, R74_61, R74_210, R74_224, R74_362, R74_386, Q74_17, Q74_61, Q74_210, Q74_224, Q74_362, Q74_386, clk );
CNU_6 CNU75(R75_18, R75_62, R75_211, R75_225, R75_363, R75_387, Q75_18, Q75_62, Q75_211, Q75_225, Q75_363, Q75_387, clk );
CNU_6 CNU76(R76_19, R76_63, R76_212, R76_226, R76_364, R76_388, Q76_19, Q76_63, Q76_212, Q76_226, Q76_364, Q76_388, clk );
CNU_6 CNU77(R77_20, R77_64, R77_213, R77_227, R77_365, R77_389, Q77_20, Q77_64, Q77_213, Q77_227, Q77_365, Q77_389, clk );
CNU_6 CNU78(R78_21, R78_65, R78_214, R78_228, R78_366, R78_390, Q78_21, Q78_65, Q78_214, Q78_228, Q78_366, Q78_390, clk );
CNU_6 CNU79(R79_22, R79_66, R79_215, R79_229, R79_367, R79_391, Q79_22, Q79_66, Q79_215, Q79_229, Q79_367, Q79_391, clk );
CNU_6 CNU80(R80_23, R80_67, R80_216, R80_230, R80_368, R80_392, Q80_23, Q80_67, Q80_216, Q80_230, Q80_368, Q80_392, clk );
CNU_6 CNU81(R81_24, R81_68, R81_193, R81_231, R81_369, R81_393, Q81_24, Q81_68, Q81_193, Q81_231, Q81_369, Q81_393, clk );
CNU_6 CNU82(R82_1, R82_69, R82_194, R82_232, R82_370, R82_394, Q82_1, Q82_69, Q82_194, Q82_232, Q82_370, Q82_394, clk );
CNU_6 CNU83(R83_2, R83_70, R83_195, R83_233, R83_371, R83_395, Q83_2, Q83_70, Q83_195, Q83_233, Q83_371, Q83_395, clk );
CNU_6 CNU84(R84_3, R84_71, R84_196, R84_234, R84_372, R84_396, Q84_3, Q84_71, Q84_196, Q84_234, Q84_372, Q84_396, clk );
CNU_6 CNU85(R85_4, R85_72, R85_197, R85_235, R85_373, R85_397, Q85_4, Q85_72, Q85_197, Q85_235, Q85_373, Q85_397, clk );
CNU_6 CNU86(R86_5, R86_49, R86_198, R86_236, R86_374, R86_398, Q86_5, Q86_49, Q86_198, Q86_236, Q86_374, Q86_398, clk );
CNU_6 CNU87(R87_6, R87_50, R87_199, R87_237, R87_375, R87_399, Q87_6, Q87_50, Q87_199, Q87_237, Q87_375, Q87_399, clk );
CNU_6 CNU88(R88_7, R88_51, R88_200, R88_238, R88_376, R88_400, Q88_7, Q88_51, Q88_200, Q88_238, Q88_376, Q88_400, clk );
CNU_6 CNU89(R89_8, R89_52, R89_201, R89_239, R89_377, R89_401, Q89_8, Q89_52, Q89_201, Q89_239, Q89_377, Q89_401, clk );
CNU_6 CNU90(R90_9, R90_53, R90_202, R90_240, R90_378, R90_402, Q90_9, Q90_53, Q90_202, Q90_240, Q90_378, Q90_402, clk );
CNU_6 CNU91(R91_10, R91_54, R91_203, R91_217, R91_379, R91_403, Q91_10, Q91_54, Q91_203, Q91_217, Q91_379, Q91_403, clk );
CNU_6 CNU92(R92_11, R92_55, R92_204, R92_218, R92_380, R92_404, Q92_11, Q92_55, Q92_204, Q92_218, Q92_380, Q92_404, clk );
CNU_6 CNU93(R93_12, R93_56, R93_205, R93_219, R93_381, R93_405, Q93_12, Q93_56, Q93_205, Q93_219, Q93_381, Q93_405, clk );
CNU_6 CNU94(R94_13, R94_57, R94_206, R94_220, R94_382, R94_406, Q94_13, Q94_57, Q94_206, Q94_220, Q94_382, Q94_406, clk );
CNU_6 CNU95(R95_14, R95_58, R95_207, R95_221, R95_383, R95_407, Q95_14, Q95_58, Q95_207, Q95_221, Q95_383, Q95_407, clk );
CNU_6 CNU96(R96_15, R96_59, R96_208, R96_222, R96_384, R96_408, Q96_15, Q96_59, Q96_208, Q96_222, Q96_384, Q96_408, clk );
CNU_6 CNU97(R97_58, R97_166, R97_227, R97_259, R97_385, R97_409, Q97_58, Q97_166, Q97_227, Q97_259, Q97_385, Q97_409, clk );
CNU_6 CNU98(R98_59, R98_167, R98_228, R98_260, R98_386, R98_410, Q98_59, Q98_167, Q98_228, Q98_260, Q98_386, Q98_410, clk );
CNU_6 CNU99(R99_60, R99_168, R99_229, R99_261, R99_387, R99_411, Q99_60, Q99_168, Q99_229, Q99_261, Q99_387, Q99_411, clk );
CNU_6 CNU100(R100_61, R100_145, R100_230, R100_262, R100_388, R100_412, Q100_61, Q100_145, Q100_230, Q100_262, Q100_388, Q100_412, clk );
CNU_6 CNU101(R101_62, R101_146, R101_231, R101_263, R101_389, R101_413, Q101_62, Q101_146, Q101_231, Q101_263, Q101_389, Q101_413, clk );
CNU_6 CNU102(R102_63, R102_147, R102_232, R102_264, R102_390, R102_414, Q102_63, Q102_147, Q102_232, Q102_264, Q102_390, Q102_414, clk );
CNU_6 CNU103(R103_64, R103_148, R103_233, R103_241, R103_391, R103_415, Q103_64, Q103_148, Q103_233, Q103_241, Q103_391, Q103_415, clk );
CNU_6 CNU104(R104_65, R104_149, R104_234, R104_242, R104_392, R104_416, Q104_65, Q104_149, Q104_234, Q104_242, Q104_392, Q104_416, clk );
CNU_6 CNU105(R105_66, R105_150, R105_235, R105_243, R105_393, R105_417, Q105_66, Q105_150, Q105_235, Q105_243, Q105_393, Q105_417, clk );
CNU_6 CNU106(R106_67, R106_151, R106_236, R106_244, R106_394, R106_418, Q106_67, Q106_151, Q106_236, Q106_244, Q106_394, Q106_418, clk );
CNU_6 CNU107(R107_68, R107_152, R107_237, R107_245, R107_395, R107_419, Q107_68, Q107_152, Q107_237, Q107_245, Q107_395, Q107_419, clk );
CNU_6 CNU108(R108_69, R108_153, R108_238, R108_246, R108_396, R108_420, Q108_69, Q108_153, Q108_238, Q108_246, Q108_396, Q108_420, clk );
CNU_6 CNU109(R109_70, R109_154, R109_239, R109_247, R109_397, R109_421, Q109_70, Q109_154, Q109_239, Q109_247, Q109_397, Q109_421, clk );
CNU_6 CNU110(R110_71, R110_155, R110_240, R110_248, R110_398, R110_422, Q110_71, Q110_155, Q110_240, Q110_248, Q110_398, Q110_422, clk );
CNU_6 CNU111(R111_72, R111_156, R111_217, R111_249, R111_399, R111_423, Q111_72, Q111_156, Q111_217, Q111_249, Q111_399, Q111_423, clk );
CNU_6 CNU112(R112_49, R112_157, R112_218, R112_250, R112_400, R112_424, Q112_49, Q112_157, Q112_218, Q112_250, Q112_400, Q112_424, clk );
CNU_6 CNU113(R113_50, R113_158, R113_219, R113_251, R113_401, R113_425, Q113_50, Q113_158, Q113_219, Q113_251, Q113_401, Q113_425, clk );
CNU_6 CNU114(R114_51, R114_159, R114_220, R114_252, R114_402, R114_426, Q114_51, Q114_159, Q114_220, Q114_252, Q114_402, Q114_426, clk );
CNU_6 CNU115(R115_52, R115_160, R115_221, R115_253, R115_403, R115_427, Q115_52, Q115_160, Q115_221, Q115_253, Q115_403, Q115_427, clk );
CNU_6 CNU116(R116_53, R116_161, R116_222, R116_254, R116_404, R116_428, Q116_53, Q116_161, Q116_222, Q116_254, Q116_404, Q116_428, clk );
CNU_6 CNU117(R117_54, R117_162, R117_223, R117_255, R117_405, R117_429, Q117_54, Q117_162, Q117_223, Q117_255, Q117_405, Q117_429, clk );
CNU_6 CNU118(R118_55, R118_163, R118_224, R118_256, R118_406, R118_430, Q118_55, Q118_163, Q118_224, Q118_256, Q118_406, Q118_430, clk );
CNU_6 CNU119(R119_56, R119_164, R119_225, R119_257, R119_407, R119_431, Q119_56, Q119_164, Q119_225, Q119_257, Q119_407, Q119_431, clk );
CNU_6 CNU120(R120_57, R120_165, R120_226, R120_258, R120_408, R120_432, Q120_57, Q120_165, Q120_226, Q120_258, Q120_408, Q120_432, clk );
CNU_7 CNU121(R121_108, R121_131, R121_189, R121_284, R121_289, R121_409, R121_433, Q121_108, Q121_131, Q121_189, Q121_284, Q121_289, Q121_409, Q121_433, clk );
CNU_7 CNU122(R122_109, R122_132, R122_190, R122_285, R122_290, R122_410, R122_434, Q122_109, Q122_132, Q122_190, Q122_285, Q122_290, Q122_410, Q122_434, clk );
CNU_7 CNU123(R123_110, R123_133, R123_191, R123_286, R123_291, R123_411, R123_435, Q123_110, Q123_133, Q123_191, Q123_286, Q123_291, Q123_411, Q123_435, clk );
CNU_7 CNU124(R124_111, R124_134, R124_192, R124_287, R124_292, R124_412, R124_436, Q124_111, Q124_134, Q124_192, Q124_287, Q124_292, Q124_412, Q124_436, clk );
CNU_7 CNU125(R125_112, R125_135, R125_169, R125_288, R125_293, R125_413, R125_437, Q125_112, Q125_135, Q125_169, Q125_288, Q125_293, Q125_413, Q125_437, clk );
CNU_7 CNU126(R126_113, R126_136, R126_170, R126_265, R126_294, R126_414, R126_438, Q126_113, Q126_136, Q126_170, Q126_265, Q126_294, Q126_414, Q126_438, clk );
CNU_7 CNU127(R127_114, R127_137, R127_171, R127_266, R127_295, R127_415, R127_439, Q127_114, Q127_137, Q127_171, Q127_266, Q127_295, Q127_415, Q127_439, clk );
CNU_7 CNU128(R128_115, R128_138, R128_172, R128_267, R128_296, R128_416, R128_440, Q128_115, Q128_138, Q128_172, Q128_267, Q128_296, Q128_416, Q128_440, clk );
CNU_7 CNU129(R129_116, R129_139, R129_173, R129_268, R129_297, R129_417, R129_441, Q129_116, Q129_139, Q129_173, Q129_268, Q129_297, Q129_417, Q129_441, clk );
CNU_7 CNU130(R130_117, R130_140, R130_174, R130_269, R130_298, R130_418, R130_442, Q130_117, Q130_140, Q130_174, Q130_269, Q130_298, Q130_418, Q130_442, clk );
CNU_7 CNU131(R131_118, R131_141, R131_175, R131_270, R131_299, R131_419, R131_443, Q131_118, Q131_141, Q131_175, Q131_270, Q131_299, Q131_419, Q131_443, clk );
CNU_7 CNU132(R132_119, R132_142, R132_176, R132_271, R132_300, R132_420, R132_444, Q132_119, Q132_142, Q132_176, Q132_271, Q132_300, Q132_420, Q132_444, clk );
CNU_7 CNU133(R133_120, R133_143, R133_177, R133_272, R133_301, R133_421, R133_445, Q133_120, Q133_143, Q133_177, Q133_272, Q133_301, Q133_421, Q133_445, clk );
CNU_7 CNU134(R134_97, R134_144, R134_178, R134_273, R134_302, R134_422, R134_446, Q134_97, Q134_144, Q134_178, Q134_273, Q134_302, Q134_422, Q134_446, clk );
CNU_7 CNU135(R135_98, R135_121, R135_179, R135_274, R135_303, R135_423, R135_447, Q135_98, Q135_121, Q135_179, Q135_274, Q135_303, Q135_423, Q135_447, clk );
CNU_7 CNU136(R136_99, R136_122, R136_180, R136_275, R136_304, R136_424, R136_448, Q136_99, Q136_122, Q136_180, Q136_275, Q136_304, Q136_424, Q136_448, clk );
CNU_7 CNU137(R137_100, R137_123, R137_181, R137_276, R137_305, R137_425, R137_449, Q137_100, Q137_123, Q137_181, Q137_276, Q137_305, Q137_425, Q137_449, clk );
CNU_7 CNU138(R138_101, R138_124, R138_182, R138_277, R138_306, R138_426, R138_450, Q138_101, Q138_124, Q138_182, Q138_277, Q138_306, Q138_426, Q138_450, clk );
CNU_7 CNU139(R139_102, R139_125, R139_183, R139_278, R139_307, R139_427, R139_451, Q139_102, Q139_125, Q139_183, Q139_278, Q139_307, Q139_427, Q139_451, clk );
CNU_7 CNU140(R140_103, R140_126, R140_184, R140_279, R140_308, R140_428, R140_452, Q140_103, Q140_126, Q140_184, Q140_279, Q140_308, Q140_428, Q140_452, clk );
CNU_7 CNU141(R141_104, R141_127, R141_185, R141_280, R141_309, R141_429, R141_453, Q141_104, Q141_127, Q141_185, Q141_280, Q141_309, Q141_429, Q141_453, clk );
CNU_7 CNU142(R142_105, R142_128, R142_186, R142_281, R142_310, R142_430, R142_454, Q142_105, Q142_128, Q142_186, Q142_281, Q142_310, Q142_430, Q142_454, clk );
CNU_7 CNU143(R143_106, R143_129, R143_187, R143_282, R143_311, R143_431, R143_455, Q143_106, Q143_129, Q143_187, Q143_282, Q143_311, Q143_431, Q143_455, clk );
CNU_7 CNU144(R144_107, R144_130, R144_188, R144_283, R144_312, R144_432, R144_456, Q144_107, Q144_130, Q144_188, Q144_283, Q144_312, Q144_432, Q144_456, clk );
CNU_6 CNU145(R145_72, R145_86, R145_220, R145_245, R145_433, R145_457, Q145_72, Q145_86, Q145_220, Q145_245, Q145_433, Q145_457, clk );
CNU_6 CNU146(R146_49, R146_87, R146_221, R146_246, R146_434, R146_458, Q146_49, Q146_87, Q146_221, Q146_246, Q146_434, Q146_458, clk );
CNU_6 CNU147(R147_50, R147_88, R147_222, R147_247, R147_435, R147_459, Q147_50, Q147_88, Q147_222, Q147_247, Q147_435, Q147_459, clk );
CNU_6 CNU148(R148_51, R148_89, R148_223, R148_248, R148_436, R148_460, Q148_51, Q148_89, Q148_223, Q148_248, Q148_436, Q148_460, clk );
CNU_6 CNU149(R149_52, R149_90, R149_224, R149_249, R149_437, R149_461, Q149_52, Q149_90, Q149_224, Q149_249, Q149_437, Q149_461, clk );
CNU_6 CNU150(R150_53, R150_91, R150_225, R150_250, R150_438, R150_462, Q150_53, Q150_91, Q150_225, Q150_250, Q150_438, Q150_462, clk );
CNU_6 CNU151(R151_54, R151_92, R151_226, R151_251, R151_439, R151_463, Q151_54, Q151_92, Q151_226, Q151_251, Q151_439, Q151_463, clk );
CNU_6 CNU152(R152_55, R152_93, R152_227, R152_252, R152_440, R152_464, Q152_55, Q152_93, Q152_227, Q152_252, Q152_440, Q152_464, clk );
CNU_6 CNU153(R153_56, R153_94, R153_228, R153_253, R153_441, R153_465, Q153_56, Q153_94, Q153_228, Q153_253, Q153_441, Q153_465, clk );
CNU_6 CNU154(R154_57, R154_95, R154_229, R154_254, R154_442, R154_466, Q154_57, Q154_95, Q154_229, Q154_254, Q154_442, Q154_466, clk );
CNU_6 CNU155(R155_58, R155_96, R155_230, R155_255, R155_443, R155_467, Q155_58, Q155_96, Q155_230, Q155_255, Q155_443, Q155_467, clk );
CNU_6 CNU156(R156_59, R156_73, R156_231, R156_256, R156_444, R156_468, Q156_59, Q156_73, Q156_231, Q156_256, Q156_444, Q156_468, clk );
CNU_6 CNU157(R157_60, R157_74, R157_232, R157_257, R157_445, R157_469, Q157_60, Q157_74, Q157_232, Q157_257, Q157_445, Q157_469, clk );
CNU_6 CNU158(R158_61, R158_75, R158_233, R158_258, R158_446, R158_470, Q158_61, Q158_75, Q158_233, Q158_258, Q158_446, Q158_470, clk );
CNU_6 CNU159(R159_62, R159_76, R159_234, R159_259, R159_447, R159_471, Q159_62, Q159_76, Q159_234, Q159_259, Q159_447, Q159_471, clk );
CNU_6 CNU160(R160_63, R160_77, R160_235, R160_260, R160_448, R160_472, Q160_63, Q160_77, Q160_235, Q160_260, Q160_448, Q160_472, clk );
CNU_6 CNU161(R161_64, R161_78, R161_236, R161_261, R161_449, R161_473, Q161_64, Q161_78, Q161_236, Q161_261, Q161_449, Q161_473, clk );
CNU_6 CNU162(R162_65, R162_79, R162_237, R162_262, R162_450, R162_474, Q162_65, Q162_79, Q162_237, Q162_262, Q162_450, Q162_474, clk );
CNU_6 CNU163(R163_66, R163_80, R163_238, R163_263, R163_451, R163_475, Q163_66, Q163_80, Q163_238, Q163_263, Q163_451, Q163_475, clk );
CNU_6 CNU164(R164_67, R164_81, R164_239, R164_264, R164_452, R164_476, Q164_67, Q164_81, Q164_239, Q164_264, Q164_452, Q164_476, clk );
CNU_6 CNU165(R165_68, R165_82, R165_240, R165_241, R165_453, R165_477, Q165_68, Q165_82, Q165_240, Q165_241, Q165_453, Q165_477, clk );
CNU_6 CNU166(R166_69, R166_83, R166_217, R166_242, R166_454, R166_478, Q166_69, Q166_83, Q166_217, Q166_242, Q166_454, Q166_478, clk );
CNU_6 CNU167(R167_70, R167_84, R167_218, R167_243, R167_455, R167_479, Q167_70, Q167_84, Q167_218, Q167_243, Q167_455, Q167_479, clk );
CNU_6 CNU168(R168_71, R168_85, R168_219, R168_244, R168_456, R168_480, Q168_71, Q168_85, Q168_219, Q168_244, Q168_456, Q168_480, clk );
CNU_6 CNU169(R169_27, R169_67, R169_145, R169_228, R169_457, R169_481, Q169_27, Q169_67, Q169_145, Q169_228, Q169_457, Q169_481, clk );
CNU_6 CNU170(R170_28, R170_68, R170_146, R170_229, R170_458, R170_482, Q170_28, Q170_68, Q170_146, Q170_229, Q170_458, Q170_482, clk );
CNU_6 CNU171(R171_29, R171_69, R171_147, R171_230, R171_459, R171_483, Q171_29, Q171_69, Q171_147, Q171_230, Q171_459, Q171_483, clk );
CNU_6 CNU172(R172_30, R172_70, R172_148, R172_231, R172_460, R172_484, Q172_30, Q172_70, Q172_148, Q172_231, Q172_460, Q172_484, clk );
CNU_6 CNU173(R173_31, R173_71, R173_149, R173_232, R173_461, R173_485, Q173_31, Q173_71, Q173_149, Q173_232, Q173_461, Q173_485, clk );
CNU_6 CNU174(R174_32, R174_72, R174_150, R174_233, R174_462, R174_486, Q174_32, Q174_72, Q174_150, Q174_233, Q174_462, Q174_486, clk );
CNU_6 CNU175(R175_33, R175_49, R175_151, R175_234, R175_463, R175_487, Q175_33, Q175_49, Q175_151, Q175_234, Q175_463, Q175_487, clk );
CNU_6 CNU176(R176_34, R176_50, R176_152, R176_235, R176_464, R176_488, Q176_34, Q176_50, Q176_152, Q176_235, Q176_464, Q176_488, clk );
CNU_6 CNU177(R177_35, R177_51, R177_153, R177_236, R177_465, R177_489, Q177_35, Q177_51, Q177_153, Q177_236, Q177_465, Q177_489, clk );
CNU_6 CNU178(R178_36, R178_52, R178_154, R178_237, R178_466, R178_490, Q178_36, Q178_52, Q178_154, Q178_237, Q178_466, Q178_490, clk );
CNU_6 CNU179(R179_37, R179_53, R179_155, R179_238, R179_467, R179_491, Q179_37, Q179_53, Q179_155, Q179_238, Q179_467, Q179_491, clk );
CNU_6 CNU180(R180_38, R180_54, R180_156, R180_239, R180_468, R180_492, Q180_38, Q180_54, Q180_156, Q180_239, Q180_468, Q180_492, clk );
CNU_6 CNU181(R181_39, R181_55, R181_157, R181_240, R181_469, R181_493, Q181_39, Q181_55, Q181_157, Q181_240, Q181_469, Q181_493, clk );
CNU_6 CNU182(R182_40, R182_56, R182_158, R182_217, R182_470, R182_494, Q182_40, Q182_56, Q182_158, Q182_217, Q182_470, Q182_494, clk );
CNU_6 CNU183(R183_41, R183_57, R183_159, R183_218, R183_471, R183_495, Q183_41, Q183_57, Q183_159, Q183_218, Q183_471, Q183_495, clk );
CNU_6 CNU184(R184_42, R184_58, R184_160, R184_219, R184_472, R184_496, Q184_42, Q184_58, Q184_160, Q184_219, Q184_472, Q184_496, clk );
CNU_6 CNU185(R185_43, R185_59, R185_161, R185_220, R185_473, R185_497, Q185_43, Q185_59, Q185_161, Q185_220, Q185_473, Q185_497, clk );
CNU_6 CNU186(R186_44, R186_60, R186_162, R186_221, R186_474, R186_498, Q186_44, Q186_60, Q186_162, Q186_221, Q186_474, Q186_498, clk );
CNU_6 CNU187(R187_45, R187_61, R187_163, R187_222, R187_475, R187_499, Q187_45, Q187_61, Q187_163, Q187_222, Q187_475, Q187_499, clk );
CNU_6 CNU188(R188_46, R188_62, R188_164, R188_223, R188_476, R188_500, Q188_46, Q188_62, Q188_164, Q188_223, Q188_476, Q188_500, clk );
CNU_6 CNU189(R189_47, R189_63, R189_165, R189_224, R189_477, R189_501, Q189_47, Q189_63, Q189_165, Q189_224, Q189_477, Q189_501, clk );
CNU_6 CNU190(R190_48, R190_64, R190_166, R190_225, R190_478, R190_502, Q190_48, Q190_64, Q190_166, Q190_225, Q190_478, Q190_502, clk );
CNU_6 CNU191(R191_25, R191_65, R191_167, R191_226, R191_479, R191_503, Q191_25, Q191_65, Q191_167, Q191_226, Q191_479, Q191_503, clk );
CNU_6 CNU192(R192_26, R192_66, R192_168, R192_227, R192_480, R192_504, Q192_26, Q192_66, Q192_168, Q192_227, Q192_480, Q192_504, clk );
CNU_7 CNU193(R193_4, R193_117, R193_127, R193_179, R193_277, R193_481, R193_505, Q193_4, Q193_117, Q193_127, Q193_179, Q193_277, Q193_481, Q193_505, clk );
CNU_7 CNU194(R194_5, R194_118, R194_128, R194_180, R194_278, R194_482, R194_506, Q194_5, Q194_118, Q194_128, Q194_180, Q194_278, Q194_482, Q194_506, clk );
CNU_7 CNU195(R195_6, R195_119, R195_129, R195_181, R195_279, R195_483, R195_507, Q195_6, Q195_119, Q195_129, Q195_181, Q195_279, Q195_483, Q195_507, clk );
CNU_7 CNU196(R196_7, R196_120, R196_130, R196_182, R196_280, R196_484, R196_508, Q196_7, Q196_120, Q196_130, Q196_182, Q196_280, Q196_484, Q196_508, clk );
CNU_7 CNU197(R197_8, R197_97, R197_131, R197_183, R197_281, R197_485, R197_509, Q197_8, Q197_97, Q197_131, Q197_183, Q197_281, Q197_485, Q197_509, clk );
CNU_7 CNU198(R198_9, R198_98, R198_132, R198_184, R198_282, R198_486, R198_510, Q198_9, Q198_98, Q198_132, Q198_184, Q198_282, Q198_486, Q198_510, clk );
CNU_7 CNU199(R199_10, R199_99, R199_133, R199_185, R199_283, R199_487, R199_511, Q199_10, Q199_99, Q199_133, Q199_185, Q199_283, Q199_487, Q199_511, clk );
CNU_7 CNU200(R200_11, R200_100, R200_134, R200_186, R200_284, R200_488, R200_512, Q200_11, Q200_100, Q200_134, Q200_186, Q200_284, Q200_488, Q200_512, clk );
CNU_7 CNU201(R201_12, R201_101, R201_135, R201_187, R201_285, R201_489, R201_513, Q201_12, Q201_101, Q201_135, Q201_187, Q201_285, Q201_489, Q201_513, clk );
CNU_7 CNU202(R202_13, R202_102, R202_136, R202_188, R202_286, R202_490, R202_514, Q202_13, Q202_102, Q202_136, Q202_188, Q202_286, Q202_490, Q202_514, clk );
CNU_7 CNU203(R203_14, R203_103, R203_137, R203_189, R203_287, R203_491, R203_515, Q203_14, Q203_103, Q203_137, Q203_189, Q203_287, Q203_491, Q203_515, clk );
CNU_7 CNU204(R204_15, R204_104, R204_138, R204_190, R204_288, R204_492, R204_516, Q204_15, Q204_104, Q204_138, Q204_190, Q204_288, Q204_492, Q204_516, clk );
CNU_7 CNU205(R205_16, R205_105, R205_139, R205_191, R205_265, R205_493, R205_517, Q205_16, Q205_105, Q205_139, Q205_191, Q205_265, Q205_493, Q205_517, clk );
CNU_7 CNU206(R206_17, R206_106, R206_140, R206_192, R206_266, R206_494, R206_518, Q206_17, Q206_106, Q206_140, Q206_192, Q206_266, Q206_494, Q206_518, clk );
CNU_7 CNU207(R207_18, R207_107, R207_141, R207_169, R207_267, R207_495, R207_519, Q207_18, Q207_107, Q207_141, Q207_169, Q207_267, Q207_495, Q207_519, clk );
CNU_7 CNU208(R208_19, R208_108, R208_142, R208_170, R208_268, R208_496, R208_520, Q208_19, Q208_108, Q208_142, Q208_170, Q208_268, Q208_496, Q208_520, clk );
CNU_7 CNU209(R209_20, R209_109, R209_143, R209_171, R209_269, R209_497, R209_521, Q209_20, Q209_109, Q209_143, Q209_171, Q209_269, Q209_497, Q209_521, clk );
CNU_7 CNU210(R210_21, R210_110, R210_144, R210_172, R210_270, R210_498, R210_522, Q210_21, Q210_110, Q210_144, Q210_172, Q210_270, Q210_498, Q210_522, clk );
CNU_7 CNU211(R211_22, R211_111, R211_121, R211_173, R211_271, R211_499, R211_523, Q211_22, Q211_111, Q211_121, Q211_173, Q211_271, Q211_499, Q211_523, clk );
CNU_7 CNU212(R212_23, R212_112, R212_122, R212_174, R212_272, R212_500, R212_524, Q212_23, Q212_112, Q212_122, Q212_174, Q212_272, Q212_500, Q212_524, clk );
CNU_7 CNU213(R213_24, R213_113, R213_123, R213_175, R213_273, R213_501, R213_525, Q213_24, Q213_113, Q213_123, Q213_175, Q213_273, Q213_501, Q213_525, clk );
CNU_7 CNU214(R214_1, R214_114, R214_124, R214_176, R214_274, R214_502, R214_526, Q214_1, Q214_114, Q214_124, Q214_176, Q214_274, Q214_502, Q214_526, clk );
CNU_7 CNU215(R215_2, R215_115, R215_125, R215_177, R215_275, R215_503, R215_527, Q215_2, Q215_115, Q215_125, Q215_177, Q215_275, Q215_503, Q215_527, clk );
CNU_7 CNU216(R216_3, R216_116, R216_126, R216_178, R216_276, R216_504, R216_528, Q216_3, Q216_116, Q216_126, Q216_178, Q216_276, Q216_504, Q216_528, clk );
CNU_6 CNU217(R217_144, R217_183, R217_258, R217_283, R217_505, R217_529, Q217_144, Q217_183, Q217_258, Q217_283, Q217_505, Q217_529, clk );
CNU_6 CNU218(R218_121, R218_184, R218_259, R218_284, R218_506, R218_530, Q218_121, Q218_184, Q218_259, Q218_284, Q218_506, Q218_530, clk );
CNU_6 CNU219(R219_122, R219_185, R219_260, R219_285, R219_507, R219_531, Q219_122, Q219_185, Q219_260, Q219_285, Q219_507, Q219_531, clk );
CNU_6 CNU220(R220_123, R220_186, R220_261, R220_286, R220_508, R220_532, Q220_123, Q220_186, Q220_261, Q220_286, Q220_508, Q220_532, clk );
CNU_6 CNU221(R221_124, R221_187, R221_262, R221_287, R221_509, R221_533, Q221_124, Q221_187, Q221_262, Q221_287, Q221_509, Q221_533, clk );
CNU_6 CNU222(R222_125, R222_188, R222_263, R222_288, R222_510, R222_534, Q222_125, Q222_188, Q222_263, Q222_288, Q222_510, Q222_534, clk );
CNU_6 CNU223(R223_126, R223_189, R223_264, R223_265, R223_511, R223_535, Q223_126, Q223_189, Q223_264, Q223_265, Q223_511, Q223_535, clk );
CNU_6 CNU224(R224_127, R224_190, R224_241, R224_266, R224_512, R224_536, Q224_127, Q224_190, Q224_241, Q224_266, Q224_512, Q224_536, clk );
CNU_6 CNU225(R225_128, R225_191, R225_242, R225_267, R225_513, R225_537, Q225_128, Q225_191, Q225_242, Q225_267, Q225_513, Q225_537, clk );
CNU_6 CNU226(R226_129, R226_192, R226_243, R226_268, R226_514, R226_538, Q226_129, Q226_192, Q226_243, Q226_268, Q226_514, Q226_538, clk );
CNU_6 CNU227(R227_130, R227_169, R227_244, R227_269, R227_515, R227_539, Q227_130, Q227_169, Q227_244, Q227_269, Q227_515, Q227_539, clk );
CNU_6 CNU228(R228_131, R228_170, R228_245, R228_270, R228_516, R228_540, Q228_131, Q228_170, Q228_245, Q228_270, Q228_516, Q228_540, clk );
CNU_6 CNU229(R229_132, R229_171, R229_246, R229_271, R229_517, R229_541, Q229_132, Q229_171, Q229_246, Q229_271, Q229_517, Q229_541, clk );
CNU_6 CNU230(R230_133, R230_172, R230_247, R230_272, R230_518, R230_542, Q230_133, Q230_172, Q230_247, Q230_272, Q230_518, Q230_542, clk );
CNU_6 CNU231(R231_134, R231_173, R231_248, R231_273, R231_519, R231_543, Q231_134, Q231_173, Q231_248, Q231_273, Q231_519, Q231_543, clk );
CNU_6 CNU232(R232_135, R232_174, R232_249, R232_274, R232_520, R232_544, Q232_135, Q232_174, Q232_249, Q232_274, Q232_520, Q232_544, clk );
CNU_6 CNU233(R233_136, R233_175, R233_250, R233_275, R233_521, R233_545, Q233_136, Q233_175, Q233_250, Q233_275, Q233_521, Q233_545, clk );
CNU_6 CNU234(R234_137, R234_176, R234_251, R234_276, R234_522, R234_546, Q234_137, Q234_176, Q234_251, Q234_276, Q234_522, Q234_546, clk );
CNU_6 CNU235(R235_138, R235_177, R235_252, R235_277, R235_523, R235_547, Q235_138, Q235_177, Q235_252, Q235_277, Q235_523, Q235_547, clk );
CNU_6 CNU236(R236_139, R236_178, R236_253, R236_278, R236_524, R236_548, Q236_139, Q236_178, Q236_253, Q236_278, Q236_524, Q236_548, clk );
CNU_6 CNU237(R237_140, R237_179, R237_254, R237_279, R237_525, R237_549, Q237_140, Q237_179, Q237_254, Q237_279, Q237_525, Q237_549, clk );
CNU_6 CNU238(R238_141, R238_180, R238_255, R238_280, R238_526, R238_550, Q238_141, Q238_180, Q238_255, Q238_280, Q238_526, Q238_550, clk );
CNU_6 CNU239(R239_142, R239_181, R239_256, R239_281, R239_527, R239_551, Q239_142, Q239_181, Q239_256, Q239_281, Q239_527, Q239_551, clk );
CNU_6 CNU240(R240_143, R240_182, R240_257, R240_282, R240_528, R240_552, Q240_143, Q240_182, Q240_257, Q240_282, Q240_528, Q240_552, clk );
CNU_6 CNU241(R241_50, R241_89, R241_202, R241_229, R241_529, R241_553, Q241_50, Q241_89, Q241_202, Q241_229, Q241_529, Q241_553, clk );
CNU_6 CNU242(R242_51, R242_90, R242_203, R242_230, R242_530, R242_554, Q242_51, Q242_90, Q242_203, Q242_230, Q242_530, Q242_554, clk );
CNU_6 CNU243(R243_52, R243_91, R243_204, R243_231, R243_531, R243_555, Q243_52, Q243_91, Q243_204, Q243_231, Q243_531, Q243_555, clk );
CNU_6 CNU244(R244_53, R244_92, R244_205, R244_232, R244_532, R244_556, Q244_53, Q244_92, Q244_205, Q244_232, Q244_532, Q244_556, clk );
CNU_6 CNU245(R245_54, R245_93, R245_206, R245_233, R245_533, R245_557, Q245_54, Q245_93, Q245_206, Q245_233, Q245_533, Q245_557, clk );
CNU_6 CNU246(R246_55, R246_94, R246_207, R246_234, R246_534, R246_558, Q246_55, Q246_94, Q246_207, Q246_234, Q246_534, Q246_558, clk );
CNU_6 CNU247(R247_56, R247_95, R247_208, R247_235, R247_535, R247_559, Q247_56, Q247_95, Q247_208, Q247_235, Q247_535, Q247_559, clk );
CNU_6 CNU248(R248_57, R248_96, R248_209, R248_236, R248_536, R248_560, Q248_57, Q248_96, Q248_209, Q248_236, Q248_536, Q248_560, clk );
CNU_6 CNU249(R249_58, R249_73, R249_210, R249_237, R249_537, R249_561, Q249_58, Q249_73, Q249_210, Q249_237, Q249_537, Q249_561, clk );
CNU_6 CNU250(R250_59, R250_74, R250_211, R250_238, R250_538, R250_562, Q250_59, Q250_74, Q250_211, Q250_238, Q250_538, Q250_562, clk );
CNU_6 CNU251(R251_60, R251_75, R251_212, R251_239, R251_539, R251_563, Q251_60, Q251_75, Q251_212, Q251_239, Q251_539, Q251_563, clk );
CNU_6 CNU252(R252_61, R252_76, R252_213, R252_240, R252_540, R252_564, Q252_61, Q252_76, Q252_213, Q252_240, Q252_540, Q252_564, clk );
CNU_6 CNU253(R253_62, R253_77, R253_214, R253_217, R253_541, R253_565, Q253_62, Q253_77, Q253_214, Q253_217, Q253_541, Q253_565, clk );
CNU_6 CNU254(R254_63, R254_78, R254_215, R254_218, R254_542, R254_566, Q254_63, Q254_78, Q254_215, Q254_218, Q254_542, Q254_566, clk );
CNU_6 CNU255(R255_64, R255_79, R255_216, R255_219, R255_543, R255_567, Q255_64, Q255_79, Q255_216, Q255_219, Q255_543, Q255_567, clk );
CNU_6 CNU256(R256_65, R256_80, R256_193, R256_220, R256_544, R256_568, Q256_65, Q256_80, Q256_193, Q256_220, Q256_544, Q256_568, clk );
CNU_6 CNU257(R257_66, R257_81, R257_194, R257_221, R257_545, R257_569, Q257_66, Q257_81, Q257_194, Q257_221, Q257_545, Q257_569, clk );
CNU_6 CNU258(R258_67, R258_82, R258_195, R258_222, R258_546, R258_570, Q258_67, Q258_82, Q258_195, Q258_222, Q258_546, Q258_570, clk );
CNU_6 CNU259(R259_68, R259_83, R259_196, R259_223, R259_547, R259_571, Q259_68, Q259_83, Q259_196, Q259_223, Q259_547, Q259_571, clk );
CNU_6 CNU260(R260_69, R260_84, R260_197, R260_224, R260_548, R260_572, Q260_69, Q260_84, Q260_197, Q260_224, Q260_548, Q260_572, clk );
CNU_6 CNU261(R261_70, R261_85, R261_198, R261_225, R261_549, R261_573, Q261_70, Q261_85, Q261_198, Q261_225, Q261_549, Q261_573, clk );
CNU_6 CNU262(R262_71, R262_86, R262_199, R262_226, R262_550, R262_574, Q262_71, Q262_86, Q262_199, Q262_226, Q262_550, Q262_574, clk );
CNU_6 CNU263(R263_72, R263_87, R263_200, R263_227, R263_551, R263_575, Q263_72, Q263_87, Q263_200, Q263_227, Q263_551, Q263_575, clk );
CNU_6 CNU264(R264_49, R264_88, R264_201, R264_228, R264_552, R264_576, Q264_49, Q264_88, Q264_201, Q264_228, Q264_552, Q264_576, clk );
CNU_6 CNU265(R265_11, R265_137, R265_179, R265_271, R265_290, R265_553, Q265_11, Q265_137, Q265_179, Q265_271, Q265_290, Q265_553, clk );
CNU_6 CNU266(R266_12, R266_138, R266_180, R266_272, R266_291, R266_554, Q266_12, Q266_138, Q266_180, Q266_272, Q266_291, Q266_554, clk );
CNU_6 CNU267(R267_13, R267_139, R267_181, R267_273, R267_292, R267_555, Q267_13, Q267_139, Q267_181, Q267_273, Q267_292, Q267_555, clk );
CNU_6 CNU268(R268_14, R268_140, R268_182, R268_274, R268_293, R268_556, Q268_14, Q268_140, Q268_182, Q268_274, Q268_293, Q268_556, clk );
CNU_6 CNU269(R269_15, R269_141, R269_183, R269_275, R269_294, R269_557, Q269_15, Q269_141, Q269_183, Q269_275, Q269_294, Q269_557, clk );
CNU_6 CNU270(R270_16, R270_142, R270_184, R270_276, R270_295, R270_558, Q270_16, Q270_142, Q270_184, Q270_276, Q270_295, Q270_558, clk );
CNU_6 CNU271(R271_17, R271_143, R271_185, R271_277, R271_296, R271_559, Q271_17, Q271_143, Q271_185, Q271_277, Q271_296, Q271_559, clk );
CNU_6 CNU272(R272_18, R272_144, R272_186, R272_278, R272_297, R272_560, Q272_18, Q272_144, Q272_186, Q272_278, Q272_297, Q272_560, clk );
CNU_6 CNU273(R273_19, R273_121, R273_187, R273_279, R273_298, R273_561, Q273_19, Q273_121, Q273_187, Q273_279, Q273_298, Q273_561, clk );
CNU_6 CNU274(R274_20, R274_122, R274_188, R274_280, R274_299, R274_562, Q274_20, Q274_122, Q274_188, Q274_280, Q274_299, Q274_562, clk );
CNU_6 CNU275(R275_21, R275_123, R275_189, R275_281, R275_300, R275_563, Q275_21, Q275_123, Q275_189, Q275_281, Q275_300, Q275_563, clk );
CNU_6 CNU276(R276_22, R276_124, R276_190, R276_282, R276_301, R276_564, Q276_22, Q276_124, Q276_190, Q276_282, Q276_301, Q276_564, clk );
CNU_6 CNU277(R277_23, R277_125, R277_191, R277_283, R277_302, R277_565, Q277_23, Q277_125, Q277_191, Q277_283, Q277_302, Q277_565, clk );
CNU_6 CNU278(R278_24, R278_126, R278_192, R278_284, R278_303, R278_566, Q278_24, Q278_126, Q278_192, Q278_284, Q278_303, Q278_566, clk );
CNU_6 CNU279(R279_1, R279_127, R279_169, R279_285, R279_304, R279_567, Q279_1, Q279_127, Q279_169, Q279_285, Q279_304, Q279_567, clk );
CNU_6 CNU280(R280_2, R280_128, R280_170, R280_286, R280_305, R280_568, Q280_2, Q280_128, Q280_170, Q280_286, Q280_305, Q280_568, clk );
CNU_6 CNU281(R281_3, R281_129, R281_171, R281_287, R281_306, R281_569, Q281_3, Q281_129, Q281_171, Q281_287, Q281_306, Q281_569, clk );
CNU_6 CNU282(R282_4, R282_130, R282_172, R282_288, R282_307, R282_570, Q282_4, Q282_130, Q282_172, Q282_288, Q282_307, Q282_570, clk );
CNU_6 CNU283(R283_5, R283_131, R283_173, R283_265, R283_308, R283_571, Q283_5, Q283_131, Q283_173, Q283_265, Q283_308, Q283_571, clk );
CNU_6 CNU284(R284_6, R284_132, R284_174, R284_266, R284_309, R284_572, Q284_6, Q284_132, Q284_174, Q284_266, Q284_309, Q284_572, clk );
CNU_6 CNU285(R285_7, R285_133, R285_175, R285_267, R285_310, R285_573, Q285_7, Q285_133, Q285_175, Q285_267, Q285_310, Q285_573, clk );
CNU_6 CNU286(R286_8, R286_134, R286_176, R286_268, R286_311, R286_574, Q286_8, Q286_134, Q286_176, Q286_268, Q286_311, Q286_574, clk );
CNU_6 CNU287(R287_9, R287_135, R287_177, R287_269, R287_312, R287_575, Q287_9, Q287_135, Q287_177, Q287_269, Q287_312, Q287_575, clk );
CNU_6 CNU288(R288_10, R288_136, R288_178, R288_270, R288_289, R288_576, Q288_10, Q288_136, Q288_178, Q288_270, Q288_289, Q288_576, clk );



VNU_3 VNU1(Q82_1, Q214_1, Q279_1, R82_1, R214_1, R279_1, L1, P1, clk ,rst);
VNU_3 VNU2(Q83_2, Q215_2, Q280_2, R83_2, R215_2, R280_2, L2, P2, clk ,rst);
VNU_3 VNU3(Q84_3, Q216_3, Q281_3, R84_3, R216_3, R281_3, L3, P3, clk ,rst);
VNU_3 VNU4(Q85_4, Q193_4, Q282_4, R85_4, R193_4, R282_4, L4, P4, clk ,rst);
VNU_3 VNU5(Q86_5, Q194_5, Q283_5, R86_5, R194_5, R283_5, L5, P5, clk ,rst);
VNU_3 VNU6(Q87_6, Q195_6, Q284_6, R87_6, R195_6, R284_6, L6, P6, clk ,rst);
VNU_3 VNU7(Q88_7, Q196_7, Q285_7, R88_7, R196_7, R285_7, L7, P7, clk ,rst);
VNU_3 VNU8(Q89_8, Q197_8, Q286_8, R89_8, R197_8, R286_8, L8, P8, clk ,rst);
VNU_3 VNU9(Q90_9, Q198_9, Q287_9, R90_9, R198_9, R287_9, L9, P9, clk ,rst);
VNU_3 VNU10(Q91_10, Q199_10, Q288_10, R91_10, R199_10, R288_10, L10, P10, clk ,rst);
VNU_3 VNU11(Q92_11, Q200_11, Q265_11, R92_11, R200_11, R265_11, L11, P11, clk ,rst);
VNU_3 VNU12(Q93_12, Q201_12, Q266_12, R93_12, R201_12, R266_12, L12, P12, clk ,rst);
VNU_3 VNU13(Q94_13, Q202_13, Q267_13, R94_13, R202_13, R267_13, L13, P13, clk ,rst);
VNU_3 VNU14(Q95_14, Q203_14, Q268_14, R95_14, R203_14, R268_14, L14, P14, clk ,rst);
VNU_3 VNU15(Q96_15, Q204_15, Q269_15, R96_15, R204_15, R269_15, L15, P15, clk ,rst);
VNU_3 VNU16(Q73_16, Q205_16, Q270_16, R73_16, R205_16, R270_16, L16, P16, clk ,rst);
VNU_3 VNU17(Q74_17, Q206_17, Q271_17, R74_17, R206_17, R271_17, L17, P17, clk ,rst);
VNU_3 VNU18(Q75_18, Q207_18, Q272_18, R75_18, R207_18, R272_18, L18, P18, clk ,rst);
VNU_3 VNU19(Q76_19, Q208_19, Q273_19, R76_19, R208_19, R273_19, L19, P19, clk ,rst);
VNU_3 VNU20(Q77_20, Q209_20, Q274_20, R77_20, R209_20, R274_20, L20, P20, clk ,rst);
VNU_3 VNU21(Q78_21, Q210_21, Q275_21, R78_21, R210_21, R275_21, L21, P21, clk ,rst);
VNU_3 VNU22(Q79_22, Q211_22, Q276_22, R79_22, R211_22, R276_22, L22, P22, clk ,rst);
VNU_3 VNU23(Q80_23, Q212_23, Q277_23, R80_23, R212_23, R277_23, L23, P23, clk ,rst);
VNU_3 VNU24(Q81_24, Q213_24, Q278_24, R81_24, R213_24, R278_24, L24, P24, clk ,rst);
VNU_3 VNU25(Q2_25, Q43_25, Q191_25, R2_25, R43_25, R191_25, L25, P25, clk ,rst);
VNU_3 VNU26(Q3_26, Q44_26, Q192_26, R3_26, R44_26, R192_26, L26, P26, clk ,rst);
VNU_3 VNU27(Q4_27, Q45_27, Q169_27, R4_27, R45_27, R169_27, L27, P27, clk ,rst);
VNU_3 VNU28(Q5_28, Q46_28, Q170_28, R5_28, R46_28, R170_28, L28, P28, clk ,rst);
VNU_3 VNU29(Q6_29, Q47_29, Q171_29, R6_29, R47_29, R171_29, L29, P29, clk ,rst);
VNU_3 VNU30(Q7_30, Q48_30, Q172_30, R7_30, R48_30, R172_30, L30, P30, clk ,rst);
VNU_3 VNU31(Q8_31, Q25_31, Q173_31, R8_31, R25_31, R173_31, L31, P31, clk ,rst);
VNU_3 VNU32(Q9_32, Q26_32, Q174_32, R9_32, R26_32, R174_32, L32, P32, clk ,rst);
VNU_3 VNU33(Q10_33, Q27_33, Q175_33, R10_33, R27_33, R175_33, L33, P33, clk ,rst);
VNU_3 VNU34(Q11_34, Q28_34, Q176_34, R11_34, R28_34, R176_34, L34, P34, clk ,rst);
VNU_3 VNU35(Q12_35, Q29_35, Q177_35, R12_35, R29_35, R177_35, L35, P35, clk ,rst);
VNU_3 VNU36(Q13_36, Q30_36, Q178_36, R13_36, R30_36, R178_36, L36, P36, clk ,rst);
VNU_3 VNU37(Q14_37, Q31_37, Q179_37, R14_37, R31_37, R179_37, L37, P37, clk ,rst);
VNU_3 VNU38(Q15_38, Q32_38, Q180_38, R15_38, R32_38, R180_38, L38, P38, clk ,rst);
VNU_3 VNU39(Q16_39, Q33_39, Q181_39, R16_39, R33_39, R181_39, L39, P39, clk ,rst);
VNU_3 VNU40(Q17_40, Q34_40, Q182_40, R17_40, R34_40, R182_40, L40, P40, clk ,rst);
VNU_3 VNU41(Q18_41, Q35_41, Q183_41, R18_41, R35_41, R183_41, L41, P41, clk ,rst);
VNU_3 VNU42(Q19_42, Q36_42, Q184_42, R19_42, R36_42, R184_42, L42, P42, clk ,rst);
VNU_3 VNU43(Q20_43, Q37_43, Q185_43, R20_43, R37_43, R185_43, L43, P43, clk ,rst);
VNU_3 VNU44(Q21_44, Q38_44, Q186_44, R21_44, R38_44, R186_44, L44, P44, clk ,rst);
VNU_3 VNU45(Q22_45, Q39_45, Q187_45, R22_45, R39_45, R187_45, L45, P45, clk ,rst);
VNU_3 VNU46(Q23_46, Q40_46, Q188_46, R23_46, R40_46, R188_46, L46, P46, clk ,rst);
VNU_3 VNU47(Q24_47, Q41_47, Q189_47, R24_47, R41_47, R189_47, L47, P47, clk ,rst);
VNU_3 VNU48(Q1_48, Q42_48, Q190_48, R1_48, R42_48, R190_48, L48, P48, clk ,rst);
VNU_6 VNU49(Q7_49, Q86_49, Q112_49, Q146_49, Q175_49, Q264_49, R7_49, R86_49, R112_49, R146_49, R175_49, R264_49, L49, P49, clk ,rst);
VNU_6 VNU50(Q8_50, Q87_50, Q113_50, Q147_50, Q176_50, Q241_50, R8_50, R87_50, R113_50, R147_50, R176_50, R241_50, L50, P50, clk ,rst);
VNU_6 VNU51(Q9_51, Q88_51, Q114_51, Q148_51, Q177_51, Q242_51, R9_51, R88_51, R114_51, R148_51, R177_51, R242_51, L51, P51, clk ,rst);
VNU_6 VNU52(Q10_52, Q89_52, Q115_52, Q149_52, Q178_52, Q243_52, R10_52, R89_52, R115_52, R149_52, R178_52, R243_52, L52, P52, clk ,rst);
VNU_6 VNU53(Q11_53, Q90_53, Q116_53, Q150_53, Q179_53, Q244_53, R11_53, R90_53, R116_53, R150_53, R179_53, R244_53, L53, P53, clk ,rst);
VNU_6 VNU54(Q12_54, Q91_54, Q117_54, Q151_54, Q180_54, Q245_54, R12_54, R91_54, R117_54, R151_54, R180_54, R245_54, L54, P54, clk ,rst);
VNU_6 VNU55(Q13_55, Q92_55, Q118_55, Q152_55, Q181_55, Q246_55, R13_55, R92_55, R118_55, R152_55, R181_55, R246_55, L55, P55, clk ,rst);
VNU_6 VNU56(Q14_56, Q93_56, Q119_56, Q153_56, Q182_56, Q247_56, R14_56, R93_56, R119_56, R153_56, R182_56, R247_56, L56, P56, clk ,rst);
VNU_6 VNU57(Q15_57, Q94_57, Q120_57, Q154_57, Q183_57, Q248_57, R15_57, R94_57, R120_57, R154_57, R183_57, R248_57, L57, P57, clk ,rst);
VNU_6 VNU58(Q16_58, Q95_58, Q97_58, Q155_58, Q184_58, Q249_58, R16_58, R95_58, R97_58, R155_58, R184_58, R249_58, L58, P58, clk ,rst);
VNU_6 VNU59(Q17_59, Q96_59, Q98_59, Q156_59, Q185_59, Q250_59, R17_59, R96_59, R98_59, R156_59, R185_59, R250_59, L59, P59, clk ,rst);
VNU_6 VNU60(Q18_60, Q73_60, Q99_60, Q157_60, Q186_60, Q251_60, R18_60, R73_60, R99_60, R157_60, R186_60, R251_60, L60, P60, clk ,rst);
VNU_6 VNU61(Q19_61, Q74_61, Q100_61, Q158_61, Q187_61, Q252_61, R19_61, R74_61, R100_61, R158_61, R187_61, R252_61, L61, P61, clk ,rst);
VNU_6 VNU62(Q20_62, Q75_62, Q101_62, Q159_62, Q188_62, Q253_62, R20_62, R75_62, R101_62, R159_62, R188_62, R253_62, L62, P62, clk ,rst);
VNU_6 VNU63(Q21_63, Q76_63, Q102_63, Q160_63, Q189_63, Q254_63, R21_63, R76_63, R102_63, R160_63, R189_63, R254_63, L63, P63, clk ,rst);
VNU_6 VNU64(Q22_64, Q77_64, Q103_64, Q161_64, Q190_64, Q255_64, R22_64, R77_64, R103_64, R161_64, R190_64, R255_64, L64, P64, clk ,rst);
VNU_6 VNU65(Q23_65, Q78_65, Q104_65, Q162_65, Q191_65, Q256_65, R23_65, R78_65, R104_65, R162_65, R191_65, R256_65, L65, P65, clk ,rst);
VNU_6 VNU66(Q24_66, Q79_66, Q105_66, Q163_66, Q192_66, Q257_66, R24_66, R79_66, R105_66, R163_66, R192_66, R257_66, L66, P66, clk ,rst);
VNU_6 VNU67(Q1_67, Q80_67, Q106_67, Q164_67, Q169_67, Q258_67, R1_67, R80_67, R106_67, R164_67, R169_67, R258_67, L67, P67, clk ,rst);
VNU_6 VNU68(Q2_68, Q81_68, Q107_68, Q165_68, Q170_68, Q259_68, R2_68, R81_68, R107_68, R165_68, R170_68, R259_68, L68, P68, clk ,rst);
VNU_6 VNU69(Q3_69, Q82_69, Q108_69, Q166_69, Q171_69, Q260_69, R3_69, R82_69, R108_69, R166_69, R171_69, R260_69, L69, P69, clk ,rst);
VNU_6 VNU70(Q4_70, Q83_70, Q109_70, Q167_70, Q172_70, Q261_70, R4_70, R83_70, R109_70, R167_70, R172_70, R261_70, L70, P70, clk ,rst);
VNU_6 VNU71(Q5_71, Q84_71, Q110_71, Q168_71, Q173_71, Q262_71, R5_71, R84_71, R110_71, R168_71, R173_71, R262_71, L71, P71, clk ,rst);
VNU_6 VNU72(Q6_72, Q85_72, Q111_72, Q145_72, Q174_72, Q263_72, R6_72, R85_72, R111_72, R145_72, R174_72, R263_72, L72, P72, clk ,rst);
VNU_3 VNU73(Q67_73, Q156_73, Q249_73, R67_73, R156_73, R249_73, L73, P73, clk ,rst);
VNU_3 VNU74(Q68_74, Q157_74, Q250_74, R68_74, R157_74, R250_74, L74, P74, clk ,rst);
VNU_3 VNU75(Q69_75, Q158_75, Q251_75, R69_75, R158_75, R251_75, L75, P75, clk ,rst);
VNU_3 VNU76(Q70_76, Q159_76, Q252_76, R70_76, R159_76, R252_76, L76, P76, clk ,rst);
VNU_3 VNU77(Q71_77, Q160_77, Q253_77, R71_77, R160_77, R253_77, L77, P77, clk ,rst);
VNU_3 VNU78(Q72_78, Q161_78, Q254_78, R72_78, R161_78, R254_78, L78, P78, clk ,rst);
VNU_3 VNU79(Q49_79, Q162_79, Q255_79, R49_79, R162_79, R255_79, L79, P79, clk ,rst);
VNU_3 VNU80(Q50_80, Q163_80, Q256_80, R50_80, R163_80, R256_80, L80, P80, clk ,rst);
VNU_3 VNU81(Q51_81, Q164_81, Q257_81, R51_81, R164_81, R257_81, L81, P81, clk ,rst);
VNU_3 VNU82(Q52_82, Q165_82, Q258_82, R52_82, R165_82, R258_82, L82, P82, clk ,rst);
VNU_3 VNU83(Q53_83, Q166_83, Q259_83, R53_83, R166_83, R259_83, L83, P83, clk ,rst);
VNU_3 VNU84(Q54_84, Q167_84, Q260_84, R54_84, R167_84, R260_84, L84, P84, clk ,rst);
VNU_3 VNU85(Q55_85, Q168_85, Q261_85, R55_85, R168_85, R261_85, L85, P85, clk ,rst);
VNU_3 VNU86(Q56_86, Q145_86, Q262_86, R56_86, R145_86, R262_86, L86, P86, clk ,rst);
VNU_3 VNU87(Q57_87, Q146_87, Q263_87, R57_87, R146_87, R263_87, L87, P87, clk ,rst);
VNU_3 VNU88(Q58_88, Q147_88, Q264_88, R58_88, R147_88, R264_88, L88, P88, clk ,rst);
VNU_3 VNU89(Q59_89, Q148_89, Q241_89, R59_89, R148_89, R241_89, L89, P89, clk ,rst);
VNU_3 VNU90(Q60_90, Q149_90, Q242_90, R60_90, R149_90, R242_90, L90, P90, clk ,rst);
VNU_3 VNU91(Q61_91, Q150_91, Q243_91, R61_91, R150_91, R243_91, L91, P91, clk ,rst);
VNU_3 VNU92(Q62_92, Q151_92, Q244_92, R62_92, R151_92, R244_92, L92, P92, clk ,rst);
VNU_3 VNU93(Q63_93, Q152_93, Q245_93, R63_93, R152_93, R245_93, L93, P93, clk ,rst);
VNU_3 VNU94(Q64_94, Q153_94, Q246_94, R64_94, R153_94, R246_94, L94, P94, clk ,rst);
VNU_3 VNU95(Q65_95, Q154_95, Q247_95, R65_95, R154_95, R247_95, L95, P95, clk ,rst);
VNU_3 VNU96(Q66_96, Q155_96, Q248_96, R66_96, R155_96, R248_96, L96, P96, clk ,rst);
VNU_3 VNU97(Q68_97, Q134_97, Q197_97, R68_97, R134_97, R197_97, L97, P97, clk ,rst);
VNU_3 VNU98(Q69_98, Q135_98, Q198_98, R69_98, R135_98, R198_98, L98, P98, clk ,rst);
VNU_3 VNU99(Q70_99, Q136_99, Q199_99, R70_99, R136_99, R199_99, L99, P99, clk ,rst);
VNU_3 VNU100(Q71_100, Q137_100, Q200_100, R71_100, R137_100, R200_100, L100, P100, clk ,rst);
VNU_3 VNU101(Q72_101, Q138_101, Q201_101, R72_101, R138_101, R201_101, L101, P101, clk ,rst);
VNU_3 VNU102(Q49_102, Q139_102, Q202_102, R49_102, R139_102, R202_102, L102, P102, clk ,rst);
VNU_3 VNU103(Q50_103, Q140_103, Q203_103, R50_103, R140_103, R203_103, L103, P103, clk ,rst);
VNU_3 VNU104(Q51_104, Q141_104, Q204_104, R51_104, R141_104, R204_104, L104, P104, clk ,rst);
VNU_3 VNU105(Q52_105, Q142_105, Q205_105, R52_105, R142_105, R205_105, L105, P105, clk ,rst);
VNU_3 VNU106(Q53_106, Q143_106, Q206_106, R53_106, R143_106, R206_106, L106, P106, clk ,rst);
VNU_3 VNU107(Q54_107, Q144_107, Q207_107, R54_107, R144_107, R207_107, L107, P107, clk ,rst);
VNU_3 VNU108(Q55_108, Q121_108, Q208_108, R55_108, R121_108, R208_108, L108, P108, clk ,rst);
VNU_3 VNU109(Q56_109, Q122_109, Q209_109, R56_109, R122_109, R209_109, L109, P109, clk ,rst);
VNU_3 VNU110(Q57_110, Q123_110, Q210_110, R57_110, R123_110, R210_110, L110, P110, clk ,rst);
VNU_3 VNU111(Q58_111, Q124_111, Q211_111, R58_111, R124_111, R211_111, L111, P111, clk ,rst);
VNU_3 VNU112(Q59_112, Q125_112, Q212_112, R59_112, R125_112, R212_112, L112, P112, clk ,rst);
VNU_3 VNU113(Q60_113, Q126_113, Q213_113, R60_113, R126_113, R213_113, L113, P113, clk ,rst);
VNU_3 VNU114(Q61_114, Q127_114, Q214_114, R61_114, R127_114, R214_114, L114, P114, clk ,rst);
VNU_3 VNU115(Q62_115, Q128_115, Q215_115, R62_115, R128_115, R215_115, L115, P115, clk ,rst);
VNU_3 VNU116(Q63_116, Q129_116, Q216_116, R63_116, R129_116, R216_116, L116, P116, clk ,rst);
VNU_3 VNU117(Q64_117, Q130_117, Q193_117, R64_117, R130_117, R193_117, L117, P117, clk ,rst);
VNU_3 VNU118(Q65_118, Q131_118, Q194_118, R65_118, R131_118, R194_118, L118, P118, clk ,rst);
VNU_3 VNU119(Q66_119, Q132_119, Q195_119, R66_119, R132_119, R195_119, L119, P119, clk ,rst);
VNU_3 VNU120(Q67_120, Q133_120, Q196_120, R67_120, R133_120, R196_120, L120, P120, clk ,rst);
VNU_6 VNU121(Q44_121, Q53_121, Q135_121, Q211_121, Q218_121, Q273_121, R44_121, R53_121, R135_121, R211_121, R218_121, R273_121, L121, P121, clk ,rst);
VNU_6 VNU122(Q45_122, Q54_122, Q136_122, Q212_122, Q219_122, Q274_122, R45_122, R54_122, R136_122, R212_122, R219_122, R274_122, L122, P122, clk ,rst);
VNU_6 VNU123(Q46_123, Q55_123, Q137_123, Q213_123, Q220_123, Q275_123, R46_123, R55_123, R137_123, R213_123, R220_123, R275_123, L123, P123, clk ,rst);
VNU_6 VNU124(Q47_124, Q56_124, Q138_124, Q214_124, Q221_124, Q276_124, R47_124, R56_124, R138_124, R214_124, R221_124, R276_124, L124, P124, clk ,rst);
VNU_6 VNU125(Q48_125, Q57_125, Q139_125, Q215_125, Q222_125, Q277_125, R48_125, R57_125, R139_125, R215_125, R222_125, R277_125, L125, P125, clk ,rst);
VNU_6 VNU126(Q25_126, Q58_126, Q140_126, Q216_126, Q223_126, Q278_126, R25_126, R58_126, R140_126, R216_126, R223_126, R278_126, L126, P126, clk ,rst);
VNU_6 VNU127(Q26_127, Q59_127, Q141_127, Q193_127, Q224_127, Q279_127, R26_127, R59_127, R141_127, R193_127, R224_127, R279_127, L127, P127, clk ,rst);
VNU_6 VNU128(Q27_128, Q60_128, Q142_128, Q194_128, Q225_128, Q280_128, R27_128, R60_128, R142_128, R194_128, R225_128, R280_128, L128, P128, clk ,rst);
VNU_6 VNU129(Q28_129, Q61_129, Q143_129, Q195_129, Q226_129, Q281_129, R28_129, R61_129, R143_129, R195_129, R226_129, R281_129, L129, P129, clk ,rst);
VNU_6 VNU130(Q29_130, Q62_130, Q144_130, Q196_130, Q227_130, Q282_130, R29_130, R62_130, R144_130, R196_130, R227_130, R282_130, L130, P130, clk ,rst);
VNU_6 VNU131(Q30_131, Q63_131, Q121_131, Q197_131, Q228_131, Q283_131, R30_131, R63_131, R121_131, R197_131, R228_131, R283_131, L131, P131, clk ,rst);
VNU_6 VNU132(Q31_132, Q64_132, Q122_132, Q198_132, Q229_132, Q284_132, R31_132, R64_132, R122_132, R198_132, R229_132, R284_132, L132, P132, clk ,rst);
VNU_6 VNU133(Q32_133, Q65_133, Q123_133, Q199_133, Q230_133, Q285_133, R32_133, R65_133, R123_133, R199_133, R230_133, R285_133, L133, P133, clk ,rst);
VNU_6 VNU134(Q33_134, Q66_134, Q124_134, Q200_134, Q231_134, Q286_134, R33_134, R66_134, R124_134, R200_134, R231_134, R286_134, L134, P134, clk ,rst);
VNU_6 VNU135(Q34_135, Q67_135, Q125_135, Q201_135, Q232_135, Q287_135, R34_135, R67_135, R125_135, R201_135, R232_135, R287_135, L135, P135, clk ,rst);
VNU_6 VNU136(Q35_136, Q68_136, Q126_136, Q202_136, Q233_136, Q288_136, R35_136, R68_136, R126_136, R202_136, R233_136, R288_136, L136, P136, clk ,rst);
VNU_6 VNU137(Q36_137, Q69_137, Q127_137, Q203_137, Q234_137, Q265_137, R36_137, R69_137, R127_137, R203_137, R234_137, R265_137, L137, P137, clk ,rst);
VNU_6 VNU138(Q37_138, Q70_138, Q128_138, Q204_138, Q235_138, Q266_138, R37_138, R70_138, R128_138, R204_138, R235_138, R266_138, L138, P138, clk ,rst);
VNU_6 VNU139(Q38_139, Q71_139, Q129_139, Q205_139, Q236_139, Q267_139, R38_139, R71_139, R129_139, R205_139, R236_139, R267_139, L139, P139, clk ,rst);
VNU_6 VNU140(Q39_140, Q72_140, Q130_140, Q206_140, Q237_140, Q268_140, R39_140, R72_140, R130_140, R206_140, R237_140, R268_140, L140, P140, clk ,rst);
VNU_6 VNU141(Q40_141, Q49_141, Q131_141, Q207_141, Q238_141, Q269_141, R40_141, R49_141, R131_141, R207_141, R238_141, R269_141, L141, P141, clk ,rst);
VNU_6 VNU142(Q41_142, Q50_142, Q132_142, Q208_142, Q239_142, Q270_142, R41_142, R50_142, R132_142, R208_142, R239_142, R270_142, L142, P142, clk ,rst);
VNU_6 VNU143(Q42_143, Q51_143, Q133_143, Q209_143, Q240_143, Q271_143, R42_143, R51_143, R133_143, R209_143, R240_143, R271_143, L143, P143, clk ,rst);
VNU_6 VNU144(Q43_144, Q52_144, Q134_144, Q210_144, Q217_144, Q272_144, R43_144, R52_144, R134_144, R210_144, R217_144, R272_144, L144, P144, clk ,rst);
VNU_3 VNU145(Q30_145, Q100_145, Q169_145, R30_145, R100_145, R169_145, L145, P145, clk ,rst);
VNU_3 VNU146(Q31_146, Q101_146, Q170_146, R31_146, R101_146, R170_146, L146, P146, clk ,rst);
VNU_3 VNU147(Q32_147, Q102_147, Q171_147, R32_147, R102_147, R171_147, L147, P147, clk ,rst);
VNU_3 VNU148(Q33_148, Q103_148, Q172_148, R33_148, R103_148, R172_148, L148, P148, clk ,rst);
VNU_3 VNU149(Q34_149, Q104_149, Q173_149, R34_149, R104_149, R173_149, L149, P149, clk ,rst);
VNU_3 VNU150(Q35_150, Q105_150, Q174_150, R35_150, R105_150, R174_150, L150, P150, clk ,rst);
VNU_3 VNU151(Q36_151, Q106_151, Q175_151, R36_151, R106_151, R175_151, L151, P151, clk ,rst);
VNU_3 VNU152(Q37_152, Q107_152, Q176_152, R37_152, R107_152, R176_152, L152, P152, clk ,rst);
VNU_3 VNU153(Q38_153, Q108_153, Q177_153, R38_153, R108_153, R177_153, L153, P153, clk ,rst);
VNU_3 VNU154(Q39_154, Q109_154, Q178_154, R39_154, R109_154, R178_154, L154, P154, clk ,rst);
VNU_3 VNU155(Q40_155, Q110_155, Q179_155, R40_155, R110_155, R179_155, L155, P155, clk ,rst);
VNU_3 VNU156(Q41_156, Q111_156, Q180_156, R41_156, R111_156, R180_156, L156, P156, clk ,rst);
VNU_3 VNU157(Q42_157, Q112_157, Q181_157, R42_157, R112_157, R181_157, L157, P157, clk ,rst);
VNU_3 VNU158(Q43_158, Q113_158, Q182_158, R43_158, R113_158, R182_158, L158, P158, clk ,rst);
VNU_3 VNU159(Q44_159, Q114_159, Q183_159, R44_159, R114_159, R183_159, L159, P159, clk ,rst);
VNU_3 VNU160(Q45_160, Q115_160, Q184_160, R45_160, R115_160, R184_160, L160, P160, clk ,rst);
VNU_3 VNU161(Q46_161, Q116_161, Q185_161, R46_161, R116_161, R185_161, L161, P161, clk ,rst);
VNU_3 VNU162(Q47_162, Q117_162, Q186_162, R47_162, R117_162, R186_162, L162, P162, clk ,rst);
VNU_3 VNU163(Q48_163, Q118_163, Q187_163, R48_163, R118_163, R187_163, L163, P163, clk ,rst);
VNU_3 VNU164(Q25_164, Q119_164, Q188_164, R25_164, R119_164, R188_164, L164, P164, clk ,rst);
VNU_3 VNU165(Q26_165, Q120_165, Q189_165, R26_165, R120_165, R189_165, L165, P165, clk ,rst);
VNU_3 VNU166(Q27_166, Q97_166, Q190_166, R27_166, R97_166, R190_166, L166, P166, clk ,rst);
VNU_3 VNU167(Q28_167, Q98_167, Q191_167, R28_167, R98_167, R191_167, L167, P167, clk ,rst);
VNU_3 VNU168(Q29_168, Q99_168, Q192_168, R29_168, R99_168, R192_168, L168, P168, clk ,rst);
VNU_6 VNU169(Q47_169, Q65_169, Q125_169, Q207_169, Q227_169, Q279_169, R47_169, R65_169, R125_169, R207_169, R227_169, R279_169, L169, P169, clk ,rst);
VNU_6 VNU170(Q48_170, Q66_170, Q126_170, Q208_170, Q228_170, Q280_170, R48_170, R66_170, R126_170, R208_170, R228_170, R280_170, L170, P170, clk ,rst);
VNU_6 VNU171(Q25_171, Q67_171, Q127_171, Q209_171, Q229_171, Q281_171, R25_171, R67_171, R127_171, R209_171, R229_171, R281_171, L171, P171, clk ,rst);
VNU_6 VNU172(Q26_172, Q68_172, Q128_172, Q210_172, Q230_172, Q282_172, R26_172, R68_172, R128_172, R210_172, R230_172, R282_172, L172, P172, clk ,rst);
VNU_6 VNU173(Q27_173, Q69_173, Q129_173, Q211_173, Q231_173, Q283_173, R27_173, R69_173, R129_173, R211_173, R231_173, R283_173, L173, P173, clk ,rst);
VNU_6 VNU174(Q28_174, Q70_174, Q130_174, Q212_174, Q232_174, Q284_174, R28_174, R70_174, R130_174, R212_174, R232_174, R284_174, L174, P174, clk ,rst);
VNU_6 VNU175(Q29_175, Q71_175, Q131_175, Q213_175, Q233_175, Q285_175, R29_175, R71_175, R131_175, R213_175, R233_175, R285_175, L175, P175, clk ,rst);
VNU_6 VNU176(Q30_176, Q72_176, Q132_176, Q214_176, Q234_176, Q286_176, R30_176, R72_176, R132_176, R214_176, R234_176, R286_176, L176, P176, clk ,rst);
VNU_6 VNU177(Q31_177, Q49_177, Q133_177, Q215_177, Q235_177, Q287_177, R31_177, R49_177, R133_177, R215_177, R235_177, R287_177, L177, P177, clk ,rst);
VNU_6 VNU178(Q32_178, Q50_178, Q134_178, Q216_178, Q236_178, Q288_178, R32_178, R50_178, R134_178, R216_178, R236_178, R288_178, L178, P178, clk ,rst);
VNU_6 VNU179(Q33_179, Q51_179, Q135_179, Q193_179, Q237_179, Q265_179, R33_179, R51_179, R135_179, R193_179, R237_179, R265_179, L179, P179, clk ,rst);
VNU_6 VNU180(Q34_180, Q52_180, Q136_180, Q194_180, Q238_180, Q266_180, R34_180, R52_180, R136_180, R194_180, R238_180, R266_180, L180, P180, clk ,rst);
VNU_6 VNU181(Q35_181, Q53_181, Q137_181, Q195_181, Q239_181, Q267_181, R35_181, R53_181, R137_181, R195_181, R239_181, R267_181, L181, P181, clk ,rst);
VNU_6 VNU182(Q36_182, Q54_182, Q138_182, Q196_182, Q240_182, Q268_182, R36_182, R54_182, R138_182, R196_182, R240_182, R268_182, L182, P182, clk ,rst);
VNU_6 VNU183(Q37_183, Q55_183, Q139_183, Q197_183, Q217_183, Q269_183, R37_183, R55_183, R139_183, R197_183, R217_183, R269_183, L183, P183, clk ,rst);
VNU_6 VNU184(Q38_184, Q56_184, Q140_184, Q198_184, Q218_184, Q270_184, R38_184, R56_184, R140_184, R198_184, R218_184, R270_184, L184, P184, clk ,rst);
VNU_6 VNU185(Q39_185, Q57_185, Q141_185, Q199_185, Q219_185, Q271_185, R39_185, R57_185, R141_185, R199_185, R219_185, R271_185, L185, P185, clk ,rst);
VNU_6 VNU186(Q40_186, Q58_186, Q142_186, Q200_186, Q220_186, Q272_186, R40_186, R58_186, R142_186, R200_186, R220_186, R272_186, L186, P186, clk ,rst);
VNU_6 VNU187(Q41_187, Q59_187, Q143_187, Q201_187, Q221_187, Q273_187, R41_187, R59_187, R143_187, R201_187, R221_187, R273_187, L187, P187, clk ,rst);
VNU_6 VNU188(Q42_188, Q60_188, Q144_188, Q202_188, Q222_188, Q274_188, R42_188, R60_188, R144_188, R202_188, R222_188, R274_188, L188, P188, clk ,rst);
VNU_6 VNU189(Q43_189, Q61_189, Q121_189, Q203_189, Q223_189, Q275_189, R43_189, R61_189, R121_189, R203_189, R223_189, R275_189, L189, P189, clk ,rst);
VNU_6 VNU190(Q44_190, Q62_190, Q122_190, Q204_190, Q224_190, Q276_190, R44_190, R62_190, R122_190, R204_190, R224_190, R276_190, L190, P190, clk ,rst);
VNU_6 VNU191(Q45_191, Q63_191, Q123_191, Q205_191, Q225_191, Q277_191, R45_191, R63_191, R123_191, R205_191, R225_191, R277_191, L191, P191, clk ,rst);
VNU_6 VNU192(Q46_192, Q64_192, Q124_192, Q206_192, Q226_192, Q278_192, R46_192, R64_192, R124_192, R206_192, R226_192, R278_192, L192, P192, clk ,rst);
VNU_3 VNU193(Q12_193, Q81_193, Q256_193, R12_193, R81_193, R256_193, L193, P193, clk ,rst);
VNU_3 VNU194(Q13_194, Q82_194, Q257_194, R13_194, R82_194, R257_194, L194, P194, clk ,rst);
VNU_3 VNU195(Q14_195, Q83_195, Q258_195, R14_195, R83_195, R258_195, L195, P195, clk ,rst);
VNU_3 VNU196(Q15_196, Q84_196, Q259_196, R15_196, R84_196, R259_196, L196, P196, clk ,rst);
VNU_3 VNU197(Q16_197, Q85_197, Q260_197, R16_197, R85_197, R260_197, L197, P197, clk ,rst);
VNU_3 VNU198(Q17_198, Q86_198, Q261_198, R17_198, R86_198, R261_198, L198, P198, clk ,rst);
VNU_3 VNU199(Q18_199, Q87_199, Q262_199, R18_199, R87_199, R262_199, L199, P199, clk ,rst);
VNU_3 VNU200(Q19_200, Q88_200, Q263_200, R19_200, R88_200, R263_200, L200, P200, clk ,rst);
VNU_3 VNU201(Q20_201, Q89_201, Q264_201, R20_201, R89_201, R264_201, L201, P201, clk ,rst);
VNU_3 VNU202(Q21_202, Q90_202, Q241_202, R21_202, R90_202, R241_202, L202, P202, clk ,rst);
VNU_3 VNU203(Q22_203, Q91_203, Q242_203, R22_203, R91_203, R242_203, L203, P203, clk ,rst);
VNU_3 VNU204(Q23_204, Q92_204, Q243_204, R23_204, R92_204, R243_204, L204, P204, clk ,rst);
VNU_3 VNU205(Q24_205, Q93_205, Q244_205, R24_205, R93_205, R244_205, L205, P205, clk ,rst);
VNU_3 VNU206(Q1_206, Q94_206, Q245_206, R1_206, R94_206, R245_206, L206, P206, clk ,rst);
VNU_3 VNU207(Q2_207, Q95_207, Q246_207, R2_207, R95_207, R246_207, L207, P207, clk ,rst);
VNU_3 VNU208(Q3_208, Q96_208, Q247_208, R3_208, R96_208, R247_208, L208, P208, clk ,rst);
VNU_3 VNU209(Q4_209, Q73_209, Q248_209, R4_209, R73_209, R248_209, L209, P209, clk ,rst);
VNU_3 VNU210(Q5_210, Q74_210, Q249_210, R5_210, R74_210, R249_210, L210, P210, clk ,rst);
VNU_3 VNU211(Q6_211, Q75_211, Q250_211, R6_211, R75_211, R250_211, L211, P211, clk ,rst);
VNU_3 VNU212(Q7_212, Q76_212, Q251_212, R7_212, R76_212, R251_212, L212, P212, clk ,rst);
VNU_3 VNU213(Q8_213, Q77_213, Q252_213, R8_213, R77_213, R252_213, L213, P213, clk ,rst);
VNU_3 VNU214(Q9_214, Q78_214, Q253_214, R9_214, R78_214, R253_214, L214, P214, clk ,rst);
VNU_3 VNU215(Q10_215, Q79_215, Q254_215, R10_215, R79_215, R254_215, L215, P215, clk ,rst);
VNU_3 VNU216(Q11_216, Q80_216, Q255_216, R11_216, R80_216, R255_216, L216, P216, clk ,rst);
VNU_6 VNU217(Q5_217, Q91_217, Q111_217, Q166_217, Q182_217, Q253_217, R5_217, R91_217, R111_217, R166_217, R182_217, R253_217, L217, P217, clk ,rst);
VNU_6 VNU218(Q6_218, Q92_218, Q112_218, Q167_218, Q183_218, Q254_218, R6_218, R92_218, R112_218, R167_218, R183_218, R254_218, L218, P218, clk ,rst);
VNU_6 VNU219(Q7_219, Q93_219, Q113_219, Q168_219, Q184_219, Q255_219, R7_219, R93_219, R113_219, R168_219, R184_219, R255_219, L219, P219, clk ,rst);
VNU_6 VNU220(Q8_220, Q94_220, Q114_220, Q145_220, Q185_220, Q256_220, R8_220, R94_220, R114_220, R145_220, R185_220, R256_220, L220, P220, clk ,rst);
VNU_6 VNU221(Q9_221, Q95_221, Q115_221, Q146_221, Q186_221, Q257_221, R9_221, R95_221, R115_221, R146_221, R186_221, R257_221, L221, P221, clk ,rst);
VNU_6 VNU222(Q10_222, Q96_222, Q116_222, Q147_222, Q187_222, Q258_222, R10_222, R96_222, R116_222, R147_222, R187_222, R258_222, L222, P222, clk ,rst);
VNU_6 VNU223(Q11_223, Q73_223, Q117_223, Q148_223, Q188_223, Q259_223, R11_223, R73_223, R117_223, R148_223, R188_223, R259_223, L223, P223, clk ,rst);
VNU_6 VNU224(Q12_224, Q74_224, Q118_224, Q149_224, Q189_224, Q260_224, R12_224, R74_224, R118_224, R149_224, R189_224, R260_224, L224, P224, clk ,rst);
VNU_6 VNU225(Q13_225, Q75_225, Q119_225, Q150_225, Q190_225, Q261_225, R13_225, R75_225, R119_225, R150_225, R190_225, R261_225, L225, P225, clk ,rst);
VNU_6 VNU226(Q14_226, Q76_226, Q120_226, Q151_226, Q191_226, Q262_226, R14_226, R76_226, R120_226, R151_226, R191_226, R262_226, L226, P226, clk ,rst);
VNU_6 VNU227(Q15_227, Q77_227, Q97_227, Q152_227, Q192_227, Q263_227, R15_227, R77_227, R97_227, R152_227, R192_227, R263_227, L227, P227, clk ,rst);
VNU_6 VNU228(Q16_228, Q78_228, Q98_228, Q153_228, Q169_228, Q264_228, R16_228, R78_228, R98_228, R153_228, R169_228, R264_228, L228, P228, clk ,rst);
VNU_6 VNU229(Q17_229, Q79_229, Q99_229, Q154_229, Q170_229, Q241_229, R17_229, R79_229, R99_229, R154_229, R170_229, R241_229, L229, P229, clk ,rst);
VNU_6 VNU230(Q18_230, Q80_230, Q100_230, Q155_230, Q171_230, Q242_230, R18_230, R80_230, R100_230, R155_230, R171_230, R242_230, L230, P230, clk ,rst);
VNU_6 VNU231(Q19_231, Q81_231, Q101_231, Q156_231, Q172_231, Q243_231, R19_231, R81_231, R101_231, R156_231, R172_231, R243_231, L231, P231, clk ,rst);
VNU_6 VNU232(Q20_232, Q82_232, Q102_232, Q157_232, Q173_232, Q244_232, R20_232, R82_232, R102_232, R157_232, R173_232, R244_232, L232, P232, clk ,rst);
VNU_6 VNU233(Q21_233, Q83_233, Q103_233, Q158_233, Q174_233, Q245_233, R21_233, R83_233, R103_233, R158_233, R174_233, R245_233, L233, P233, clk ,rst);
VNU_6 VNU234(Q22_234, Q84_234, Q104_234, Q159_234, Q175_234, Q246_234, R22_234, R84_234, R104_234, R159_234, R175_234, R246_234, L234, P234, clk ,rst);
VNU_6 VNU235(Q23_235, Q85_235, Q105_235, Q160_235, Q176_235, Q247_235, R23_235, R85_235, R105_235, R160_235, R176_235, R247_235, L235, P235, clk ,rst);
VNU_6 VNU236(Q24_236, Q86_236, Q106_236, Q161_236, Q177_236, Q248_236, R24_236, R86_236, R106_236, R161_236, R177_236, R248_236, L236, P236, clk ,rst);
VNU_6 VNU237(Q1_237, Q87_237, Q107_237, Q162_237, Q178_237, Q249_237, R1_237, R87_237, R107_237, R162_237, R178_237, R249_237, L237, P237, clk ,rst);
VNU_6 VNU238(Q2_238, Q88_238, Q108_238, Q163_238, Q179_238, Q250_238, R2_238, R88_238, R108_238, R163_238, R179_238, R250_238, L238, P238, clk ,rst);
VNU_6 VNU239(Q3_239, Q89_239, Q109_239, Q164_239, Q180_239, Q251_239, R3_239, R89_239, R109_239, R164_239, R180_239, R251_239, L239, P239, clk ,rst);
VNU_6 VNU240(Q4_240, Q90_240, Q110_240, Q165_240, Q181_240, Q252_240, R4_240, R90_240, R110_240, R165_240, R181_240, R252_240, L240, P240, clk ,rst);
VNU_3 VNU241(Q103_241, Q165_241, Q224_241, R103_241, R165_241, R224_241, L241, P241, clk ,rst);
VNU_3 VNU242(Q104_242, Q166_242, Q225_242, R104_242, R166_242, R225_242, L242, P242, clk ,rst);
VNU_3 VNU243(Q105_243, Q167_243, Q226_243, R105_243, R167_243, R226_243, L243, P243, clk ,rst);
VNU_3 VNU244(Q106_244, Q168_244, Q227_244, R106_244, R168_244, R227_244, L244, P244, clk ,rst);
VNU_3 VNU245(Q107_245, Q145_245, Q228_245, R107_245, R145_245, R228_245, L245, P245, clk ,rst);
VNU_3 VNU246(Q108_246, Q146_246, Q229_246, R108_246, R146_246, R229_246, L246, P246, clk ,rst);
VNU_3 VNU247(Q109_247, Q147_247, Q230_247, R109_247, R147_247, R230_247, L247, P247, clk ,rst);
VNU_3 VNU248(Q110_248, Q148_248, Q231_248, R110_248, R148_248, R231_248, L248, P248, clk ,rst);
VNU_3 VNU249(Q111_249, Q149_249, Q232_249, R111_249, R149_249, R232_249, L249, P249, clk ,rst);
VNU_3 VNU250(Q112_250, Q150_250, Q233_250, R112_250, R150_250, R233_250, L250, P250, clk ,rst);
VNU_3 VNU251(Q113_251, Q151_251, Q234_251, R113_251, R151_251, R234_251, L251, P251, clk ,rst);
VNU_3 VNU252(Q114_252, Q152_252, Q235_252, R114_252, R152_252, R235_252, L252, P252, clk ,rst);
VNU_3 VNU253(Q115_253, Q153_253, Q236_253, R115_253, R153_253, R236_253, L253, P253, clk ,rst);
VNU_3 VNU254(Q116_254, Q154_254, Q237_254, R116_254, R154_254, R237_254, L254, P254, clk ,rst);
VNU_3 VNU255(Q117_255, Q155_255, Q238_255, R117_255, R155_255, R238_255, L255, P255, clk ,rst);
VNU_3 VNU256(Q118_256, Q156_256, Q239_256, R118_256, R156_256, R239_256, L256, P256, clk ,rst);
VNU_3 VNU257(Q119_257, Q157_257, Q240_257, R119_257, R157_257, R240_257, L257, P257, clk ,rst);
VNU_3 VNU258(Q120_258, Q158_258, Q217_258, R120_258, R158_258, R217_258, L258, P258, clk ,rst);
VNU_3 VNU259(Q97_259, Q159_259, Q218_259, R97_259, R159_259, R218_259, L259, P259, clk ,rst);
VNU_3 VNU260(Q98_260, Q160_260, Q219_260, R98_260, R160_260, R219_260, L260, P260, clk ,rst);
VNU_3 VNU261(Q99_261, Q161_261, Q220_261, R99_261, R161_261, R220_261, L261, P261, clk ,rst);
VNU_3 VNU262(Q100_262, Q162_262, Q221_262, R100_262, R162_262, R221_262, L262, P262, clk ,rst);
VNU_3 VNU263(Q101_263, Q163_263, Q222_263, R101_263, R163_263, R222_263, L263, P263, clk ,rst);
VNU_3 VNU264(Q102_264, Q164_264, Q223_264, R102_264, R164_264, R223_264, L264, P264, clk ,rst);
VNU_6 VNU265(Q46_265, Q49_265, Q126_265, Q205_265, Q223_265, Q283_265, R46_265, R49_265, R126_265, R205_265, R223_265, R283_265, L265, P265, clk ,rst);
VNU_6 VNU266(Q47_266, Q50_266, Q127_266, Q206_266, Q224_266, Q284_266, R47_266, R50_266, R127_266, R206_266, R224_266, R284_266, L266, P266, clk ,rst);
VNU_6 VNU267(Q48_267, Q51_267, Q128_267, Q207_267, Q225_267, Q285_267, R48_267, R51_267, R128_267, R207_267, R225_267, R285_267, L267, P267, clk ,rst);
VNU_6 VNU268(Q25_268, Q52_268, Q129_268, Q208_268, Q226_268, Q286_268, R25_268, R52_268, R129_268, R208_268, R226_268, R286_268, L268, P268, clk ,rst);
VNU_6 VNU269(Q26_269, Q53_269, Q130_269, Q209_269, Q227_269, Q287_269, R26_269, R53_269, R130_269, R209_269, R227_269, R287_269, L269, P269, clk ,rst);
VNU_6 VNU270(Q27_270, Q54_270, Q131_270, Q210_270, Q228_270, Q288_270, R27_270, R54_270, R131_270, R210_270, R228_270, R288_270, L270, P270, clk ,rst);
VNU_6 VNU271(Q28_271, Q55_271, Q132_271, Q211_271, Q229_271, Q265_271, R28_271, R55_271, R132_271, R211_271, R229_271, R265_271, L271, P271, clk ,rst);
VNU_6 VNU272(Q29_272, Q56_272, Q133_272, Q212_272, Q230_272, Q266_272, R29_272, R56_272, R133_272, R212_272, R230_272, R266_272, L272, P272, clk ,rst);
VNU_6 VNU273(Q30_273, Q57_273, Q134_273, Q213_273, Q231_273, Q267_273, R30_273, R57_273, R134_273, R213_273, R231_273, R267_273, L273, P273, clk ,rst);
VNU_6 VNU274(Q31_274, Q58_274, Q135_274, Q214_274, Q232_274, Q268_274, R31_274, R58_274, R135_274, R214_274, R232_274, R268_274, L274, P274, clk ,rst);
VNU_6 VNU275(Q32_275, Q59_275, Q136_275, Q215_275, Q233_275, Q269_275, R32_275, R59_275, R136_275, R215_275, R233_275, R269_275, L275, P275, clk ,rst);
VNU_6 VNU276(Q33_276, Q60_276, Q137_276, Q216_276, Q234_276, Q270_276, R33_276, R60_276, R137_276, R216_276, R234_276, R270_276, L276, P276, clk ,rst);
VNU_6 VNU277(Q34_277, Q61_277, Q138_277, Q193_277, Q235_277, Q271_277, R34_277, R61_277, R138_277, R193_277, R235_277, R271_277, L277, P277, clk ,rst);
VNU_6 VNU278(Q35_278, Q62_278, Q139_278, Q194_278, Q236_278, Q272_278, R35_278, R62_278, R139_278, R194_278, R236_278, R272_278, L278, P278, clk ,rst);
VNU_6 VNU279(Q36_279, Q63_279, Q140_279, Q195_279, Q237_279, Q273_279, R36_279, R63_279, R140_279, R195_279, R237_279, R273_279, L279, P279, clk ,rst);
VNU_6 VNU280(Q37_280, Q64_280, Q141_280, Q196_280, Q238_280, Q274_280, R37_280, R64_280, R141_280, R196_280, R238_280, R274_280, L280, P280, clk ,rst);
VNU_6 VNU281(Q38_281, Q65_281, Q142_281, Q197_281, Q239_281, Q275_281, R38_281, R65_281, R142_281, R197_281, R239_281, R275_281, L281, P281, clk ,rst);
VNU_6 VNU282(Q39_282, Q66_282, Q143_282, Q198_282, Q240_282, Q276_282, R39_282, R66_282, R143_282, R198_282, R240_282, R276_282, L282, P282, clk ,rst);
VNU_6 VNU283(Q40_283, Q67_283, Q144_283, Q199_283, Q217_283, Q277_283, R40_283, R67_283, R144_283, R199_283, R217_283, R277_283, L283, P283, clk ,rst);
VNU_6 VNU284(Q41_284, Q68_284, Q121_284, Q200_284, Q218_284, Q278_284, R41_284, R68_284, R121_284, R200_284, R218_284, R278_284, L284, P284, clk ,rst);
VNU_6 VNU285(Q42_285, Q69_285, Q122_285, Q201_285, Q219_285, Q279_285, R42_285, R69_285, R122_285, R201_285, R219_285, R279_285, L285, P285, clk ,rst);
VNU_6 VNU286(Q43_286, Q70_286, Q123_286, Q202_286, Q220_286, Q280_286, R43_286, R70_286, R123_286, R202_286, R220_286, R280_286, L286, P286, clk ,rst);
VNU_6 VNU287(Q44_287, Q71_287, Q124_287, Q203_287, Q221_287, Q281_287, R44_287, R71_287, R124_287, R203_287, R221_287, R281_287, L287, P287, clk ,rst);
VNU_6 VNU288(Q45_288, Q72_288, Q125_288, Q204_288, Q222_288, Q282_288, R45_288, R72_288, R125_288, R204_288, R222_288, R282_288, L288, P288, clk ,rst);
VNU_3 VNU289(Q24_289, Q121_289, Q288_289, R24_289, R121_289, R288_289, L289, P289, clk ,rst);
VNU_3 VNU290(Q1_290, Q122_290, Q265_290, R1_290, R122_290, R265_290, L290, P290, clk ,rst);
VNU_3 VNU291(Q2_291, Q123_291, Q266_291, R2_291, R123_291, R266_291, L291, P291, clk ,rst);
VNU_3 VNU292(Q3_292, Q124_292, Q267_292, R3_292, R124_292, R267_292, L292, P292, clk ,rst);
VNU_3 VNU293(Q4_293, Q125_293, Q268_293, R4_293, R125_293, R268_293, L293, P293, clk ,rst);
VNU_3 VNU294(Q5_294, Q126_294, Q269_294, R5_294, R126_294, R269_294, L294, P294, clk ,rst);
VNU_3 VNU295(Q6_295, Q127_295, Q270_295, R6_295, R127_295, R270_295, L295, P295, clk ,rst);
VNU_3 VNU296(Q7_296, Q128_296, Q271_296, R7_296, R128_296, R271_296, L296, P296, clk ,rst);
VNU_3 VNU297(Q8_297, Q129_297, Q272_297, R8_297, R129_297, R272_297, L297, P297, clk ,rst);
VNU_3 VNU298(Q9_298, Q130_298, Q273_298, R9_298, R130_298, R273_298, L298, P298, clk ,rst);
VNU_3 VNU299(Q10_299, Q131_299, Q274_299, R10_299, R131_299, R274_299, L299, P299, clk ,rst);
VNU_3 VNU300(Q11_300, Q132_300, Q275_300, R11_300, R132_300, R275_300, L300, P300, clk ,rst);
VNU_3 VNU301(Q12_301, Q133_301, Q276_301, R12_301, R133_301, R276_301, L301, P301, clk ,rst);
VNU_3 VNU302(Q13_302, Q134_302, Q277_302, R13_302, R134_302, R277_302, L302, P302, clk ,rst);
VNU_3 VNU303(Q14_303, Q135_303, Q278_303, R14_303, R135_303, R278_303, L303, P303, clk ,rst);
VNU_3 VNU304(Q15_304, Q136_304, Q279_304, R15_304, R136_304, R279_304, L304, P304, clk ,rst);
VNU_3 VNU305(Q16_305, Q137_305, Q280_305, R16_305, R137_305, R280_305, L305, P305, clk ,rst);
VNU_3 VNU306(Q17_306, Q138_306, Q281_306, R17_306, R138_306, R281_306, L306, P306, clk ,rst);
VNU_3 VNU307(Q18_307, Q139_307, Q282_307, R18_307, R139_307, R282_307, L307, P307, clk ,rst);
VNU_3 VNU308(Q19_308, Q140_308, Q283_308, R19_308, R140_308, R283_308, L308, P308, clk ,rst);
VNU_3 VNU309(Q20_309, Q141_309, Q284_309, R20_309, R141_309, R284_309, L309, P309, clk ,rst);
VNU_3 VNU310(Q21_310, Q142_310, Q285_310, R21_310, R142_310, R285_310, L310, P310, clk ,rst);
VNU_3 VNU311(Q22_311, Q143_311, Q286_311, R22_311, R143_311, R286_311, L311, P311, clk ,rst);
VNU_3 VNU312(Q23_312, Q144_312, Q287_312, R23_312, R144_312, R287_312, L312, P312, clk ,rst);
VNU_2 VNU313(Q1_313, Q25_313, R1_313, R25_313, L313, P313, clk ,rst);
VNU_2 VNU314(Q2_314, Q26_314, R2_314, R26_314, L314, P314, clk ,rst);
VNU_2 VNU315(Q3_315, Q27_315, R3_315, R27_315, L315, P315, clk ,rst);
VNU_2 VNU316(Q4_316, Q28_316, R4_316, R28_316, L316, P316, clk ,rst);
VNU_2 VNU317(Q5_317, Q29_317, R5_317, R29_317, L317, P317, clk ,rst);
VNU_2 VNU318(Q6_318, Q30_318, R6_318, R30_318, L318, P318, clk ,rst);
VNU_2 VNU319(Q7_319, Q31_319, R7_319, R31_319, L319, P319, clk ,rst);
VNU_2 VNU320(Q8_320, Q32_320, R8_320, R32_320, L320, P320, clk ,rst);
VNU_2 VNU321(Q9_321, Q33_321, R9_321, R33_321, L321, P321, clk ,rst);
VNU_2 VNU322(Q10_322, Q34_322, R10_322, R34_322, L322, P322, clk ,rst);
VNU_2 VNU323(Q11_323, Q35_323, R11_323, R35_323, L323, P323, clk ,rst);
VNU_2 VNU324(Q12_324, Q36_324, R12_324, R36_324, L324, P324, clk ,rst);
VNU_2 VNU325(Q13_325, Q37_325, R13_325, R37_325, L325, P325, clk ,rst);
VNU_2 VNU326(Q14_326, Q38_326, R14_326, R38_326, L326, P326, clk ,rst);
VNU_2 VNU327(Q15_327, Q39_327, R15_327, R39_327, L327, P327, clk ,rst);
VNU_2 VNU328(Q16_328, Q40_328, R16_328, R40_328, L328, P328, clk ,rst);
VNU_2 VNU329(Q17_329, Q41_329, R17_329, R41_329, L329, P329, clk ,rst);
VNU_2 VNU330(Q18_330, Q42_330, R18_330, R42_330, L330, P330, clk ,rst);
VNU_2 VNU331(Q19_331, Q43_331, R19_331, R43_331, L331, P331, clk ,rst);
VNU_2 VNU332(Q20_332, Q44_332, R20_332, R44_332, L332, P332, clk ,rst);
VNU_2 VNU333(Q21_333, Q45_333, R21_333, R45_333, L333, P333, clk ,rst);
VNU_2 VNU334(Q22_334, Q46_334, R22_334, R46_334, L334, P334, clk ,rst);
VNU_2 VNU335(Q23_335, Q47_335, R23_335, R47_335, L335, P335, clk ,rst);
VNU_2 VNU336(Q24_336, Q48_336, R24_336, R48_336, L336, P336, clk ,rst);
VNU_2 VNU337(Q25_337, Q49_337, R25_337, R49_337, L337, P337, clk ,rst);
VNU_2 VNU338(Q26_338, Q50_338, R26_338, R50_338, L338, P338, clk ,rst);
VNU_2 VNU339(Q27_339, Q51_339, R27_339, R51_339, L339, P339, clk ,rst);
VNU_2 VNU340(Q28_340, Q52_340, R28_340, R52_340, L340, P340, clk ,rst);
VNU_2 VNU341(Q29_341, Q53_341, R29_341, R53_341, L341, P341, clk ,rst);
VNU_2 VNU342(Q30_342, Q54_342, R30_342, R54_342, L342, P342, clk ,rst);
VNU_2 VNU343(Q31_343, Q55_343, R31_343, R55_343, L343, P343, clk ,rst);
VNU_2 VNU344(Q32_344, Q56_344, R32_344, R56_344, L344, P344, clk ,rst);
VNU_2 VNU345(Q33_345, Q57_345, R33_345, R57_345, L345, P345, clk ,rst);
VNU_2 VNU346(Q34_346, Q58_346, R34_346, R58_346, L346, P346, clk ,rst);
VNU_2 VNU347(Q35_347, Q59_347, R35_347, R59_347, L347, P347, clk ,rst);
VNU_2 VNU348(Q36_348, Q60_348, R36_348, R60_348, L348, P348, clk ,rst);
VNU_2 VNU349(Q37_349, Q61_349, R37_349, R61_349, L349, P349, clk ,rst);
VNU_2 VNU350(Q38_350, Q62_350, R38_350, R62_350, L350, P350, clk ,rst);
VNU_2 VNU351(Q39_351, Q63_351, R39_351, R63_351, L351, P351, clk ,rst);
VNU_2 VNU352(Q40_352, Q64_352, R40_352, R64_352, L352, P352, clk ,rst);
VNU_2 VNU353(Q41_353, Q65_353, R41_353, R65_353, L353, P353, clk ,rst);
VNU_2 VNU354(Q42_354, Q66_354, R42_354, R66_354, L354, P354, clk ,rst);
VNU_2 VNU355(Q43_355, Q67_355, R43_355, R67_355, L355, P355, clk ,rst);
VNU_2 VNU356(Q44_356, Q68_356, R44_356, R68_356, L356, P356, clk ,rst);
VNU_2 VNU357(Q45_357, Q69_357, R45_357, R69_357, L357, P357, clk ,rst);
VNU_2 VNU358(Q46_358, Q70_358, R46_358, R70_358, L358, P358, clk ,rst);
VNU_2 VNU359(Q47_359, Q71_359, R47_359, R71_359, L359, P359, clk ,rst);
VNU_2 VNU360(Q48_360, Q72_360, R48_360, R72_360, L360, P360, clk ,rst);
VNU_2 VNU361(Q49_361, Q73_361, R49_361, R73_361, L361, P361, clk ,rst);
VNU_2 VNU362(Q50_362, Q74_362, R50_362, R74_362, L362, P362, clk ,rst);
VNU_2 VNU363(Q51_363, Q75_363, R51_363, R75_363, L363, P363, clk ,rst);
VNU_2 VNU364(Q52_364, Q76_364, R52_364, R76_364, L364, P364, clk ,rst);
VNU_2 VNU365(Q53_365, Q77_365, R53_365, R77_365, L365, P365, clk ,rst);
VNU_2 VNU366(Q54_366, Q78_366, R54_366, R78_366, L366, P366, clk ,rst);
VNU_2 VNU367(Q55_367, Q79_367, R55_367, R79_367, L367, P367, clk ,rst);
VNU_2 VNU368(Q56_368, Q80_368, R56_368, R80_368, L368, P368, clk ,rst);
VNU_2 VNU369(Q57_369, Q81_369, R57_369, R81_369, L369, P369, clk ,rst);
VNU_2 VNU370(Q58_370, Q82_370, R58_370, R82_370, L370, P370, clk ,rst);
VNU_2 VNU371(Q59_371, Q83_371, R59_371, R83_371, L371, P371, clk ,rst);
VNU_2 VNU372(Q60_372, Q84_372, R60_372, R84_372, L372, P372, clk ,rst);
VNU_2 VNU373(Q61_373, Q85_373, R61_373, R85_373, L373, P373, clk ,rst);
VNU_2 VNU374(Q62_374, Q86_374, R62_374, R86_374, L374, P374, clk ,rst);
VNU_2 VNU375(Q63_375, Q87_375, R63_375, R87_375, L375, P375, clk ,rst);
VNU_2 VNU376(Q64_376, Q88_376, R64_376, R88_376, L376, P376, clk ,rst);
VNU_2 VNU377(Q65_377, Q89_377, R65_377, R89_377, L377, P377, clk ,rst);
VNU_2 VNU378(Q66_378, Q90_378, R66_378, R90_378, L378, P378, clk ,rst);
VNU_2 VNU379(Q67_379, Q91_379, R67_379, R91_379, L379, P379, clk ,rst);
VNU_2 VNU380(Q68_380, Q92_380, R68_380, R92_380, L380, P380, clk ,rst);
VNU_2 VNU381(Q69_381, Q93_381, R69_381, R93_381, L381, P381, clk ,rst);
VNU_2 VNU382(Q70_382, Q94_382, R70_382, R94_382, L382, P382, clk ,rst);
VNU_2 VNU383(Q71_383, Q95_383, R71_383, R95_383, L383, P383, clk ,rst);
VNU_2 VNU384(Q72_384, Q96_384, R72_384, R96_384, L384, P384, clk ,rst);
VNU_2 VNU385(Q73_385, Q97_385, R73_385, R97_385, L385, P385, clk ,rst);
VNU_2 VNU386(Q74_386, Q98_386, R74_386, R98_386, L386, P386, clk ,rst);
VNU_2 VNU387(Q75_387, Q99_387, R75_387, R99_387, L387, P387, clk ,rst);
VNU_2 VNU388(Q76_388, Q100_388, R76_388, R100_388, L388, P388, clk ,rst);
VNU_2 VNU389(Q77_389, Q101_389, R77_389, R101_389, L389, P389, clk ,rst);
VNU_2 VNU390(Q78_390, Q102_390, R78_390, R102_390, L390, P390, clk ,rst);
VNU_2 VNU391(Q79_391, Q103_391, R79_391, R103_391, L391, P391, clk ,rst);
VNU_2 VNU392(Q80_392, Q104_392, R80_392, R104_392, L392, P392, clk ,rst);
VNU_2 VNU393(Q81_393, Q105_393, R81_393, R105_393, L393, P393, clk ,rst);
VNU_2 VNU394(Q82_394, Q106_394, R82_394, R106_394, L394, P394, clk ,rst);
VNU_2 VNU395(Q83_395, Q107_395, R83_395, R107_395, L395, P395, clk ,rst);
VNU_2 VNU396(Q84_396, Q108_396, R84_396, R108_396, L396, P396, clk ,rst);
VNU_2 VNU397(Q85_397, Q109_397, R85_397, R109_397, L397, P397, clk ,rst);
VNU_2 VNU398(Q86_398, Q110_398, R86_398, R110_398, L398, P398, clk ,rst);
VNU_2 VNU399(Q87_399, Q111_399, R87_399, R111_399, L399, P399, clk ,rst);
VNU_2 VNU400(Q88_400, Q112_400, R88_400, R112_400, L400, P400, clk ,rst);
VNU_2 VNU401(Q89_401, Q113_401, R89_401, R113_401, L401, P401, clk ,rst);
VNU_2 VNU402(Q90_402, Q114_402, R90_402, R114_402, L402, P402, clk ,rst);
VNU_2 VNU403(Q91_403, Q115_403, R91_403, R115_403, L403, P403, clk ,rst);
VNU_2 VNU404(Q92_404, Q116_404, R92_404, R116_404, L404, P404, clk ,rst);
VNU_2 VNU405(Q93_405, Q117_405, R93_405, R117_405, L405, P405, clk ,rst);
VNU_2 VNU406(Q94_406, Q118_406, R94_406, R118_406, L406, P406, clk ,rst);
VNU_2 VNU407(Q95_407, Q119_407, R95_407, R119_407, L407, P407, clk ,rst);
VNU_2 VNU408(Q96_408, Q120_408, R96_408, R120_408, L408, P408, clk ,rst);
VNU_2 VNU409(Q97_409, Q121_409, R97_409, R121_409, L409, P409, clk ,rst);
VNU_2 VNU410(Q98_410, Q122_410, R98_410, R122_410, L410, P410, clk ,rst);
VNU_2 VNU411(Q99_411, Q123_411, R99_411, R123_411, L411, P411, clk ,rst);
VNU_2 VNU412(Q100_412, Q124_412, R100_412, R124_412, L412, P412, clk ,rst);
VNU_2 VNU413(Q101_413, Q125_413, R101_413, R125_413, L413, P413, clk ,rst);
VNU_2 VNU414(Q102_414, Q126_414, R102_414, R126_414, L414, P414, clk ,rst);
VNU_2 VNU415(Q103_415, Q127_415, R103_415, R127_415, L415, P415, clk ,rst);
VNU_2 VNU416(Q104_416, Q128_416, R104_416, R128_416, L416, P416, clk ,rst);
VNU_2 VNU417(Q105_417, Q129_417, R105_417, R129_417, L417, P417, clk ,rst);
VNU_2 VNU418(Q106_418, Q130_418, R106_418, R130_418, L418, P418, clk ,rst);
VNU_2 VNU419(Q107_419, Q131_419, R107_419, R131_419, L419, P419, clk ,rst);
VNU_2 VNU420(Q108_420, Q132_420, R108_420, R132_420, L420, P420, clk ,rst);
VNU_2 VNU421(Q109_421, Q133_421, R109_421, R133_421, L421, P421, clk ,rst);
VNU_2 VNU422(Q110_422, Q134_422, R110_422, R134_422, L422, P422, clk ,rst);
VNU_2 VNU423(Q111_423, Q135_423, R111_423, R135_423, L423, P423, clk ,rst);
VNU_2 VNU424(Q112_424, Q136_424, R112_424, R136_424, L424, P424, clk ,rst);
VNU_2 VNU425(Q113_425, Q137_425, R113_425, R137_425, L425, P425, clk ,rst);
VNU_2 VNU426(Q114_426, Q138_426, R114_426, R138_426, L426, P426, clk ,rst);
VNU_2 VNU427(Q115_427, Q139_427, R115_427, R139_427, L427, P427, clk ,rst);
VNU_2 VNU428(Q116_428, Q140_428, R116_428, R140_428, L428, P428, clk ,rst);
VNU_2 VNU429(Q117_429, Q141_429, R117_429, R141_429, L429, P429, clk ,rst);
VNU_2 VNU430(Q118_430, Q142_430, R118_430, R142_430, L430, P430, clk ,rst);
VNU_2 VNU431(Q119_431, Q143_431, R119_431, R143_431, L431, P431, clk ,rst);
VNU_2 VNU432(Q120_432, Q144_432, R120_432, R144_432, L432, P432, clk ,rst);
VNU_2 VNU433(Q121_433, Q145_433, R121_433, R145_433, L433, P433, clk ,rst);
VNU_2 VNU434(Q122_434, Q146_434, R122_434, R146_434, L434, P434, clk ,rst);
VNU_2 VNU435(Q123_435, Q147_435, R123_435, R147_435, L435, P435, clk ,rst);
VNU_2 VNU436(Q124_436, Q148_436, R124_436, R148_436, L436, P436, clk ,rst);
VNU_2 VNU437(Q125_437, Q149_437, R125_437, R149_437, L437, P437, clk ,rst);
VNU_2 VNU438(Q126_438, Q150_438, R126_438, R150_438, L438, P438, clk ,rst);
VNU_2 VNU439(Q127_439, Q151_439, R127_439, R151_439, L439, P439, clk ,rst);
VNU_2 VNU440(Q128_440, Q152_440, R128_440, R152_440, L440, P440, clk ,rst);
VNU_2 VNU441(Q129_441, Q153_441, R129_441, R153_441, L441, P441, clk ,rst);
VNU_2 VNU442(Q130_442, Q154_442, R130_442, R154_442, L442, P442, clk ,rst);
VNU_2 VNU443(Q131_443, Q155_443, R131_443, R155_443, L443, P443, clk ,rst);
VNU_2 VNU444(Q132_444, Q156_444, R132_444, R156_444, L444, P444, clk ,rst);
VNU_2 VNU445(Q133_445, Q157_445, R133_445, R157_445, L445, P445, clk ,rst);
VNU_2 VNU446(Q134_446, Q158_446, R134_446, R158_446, L446, P446, clk ,rst);
VNU_2 VNU447(Q135_447, Q159_447, R135_447, R159_447, L447, P447, clk ,rst);
VNU_2 VNU448(Q136_448, Q160_448, R136_448, R160_448, L448, P448, clk ,rst);
VNU_2 VNU449(Q137_449, Q161_449, R137_449, R161_449, L449, P449, clk ,rst);
VNU_2 VNU450(Q138_450, Q162_450, R138_450, R162_450, L450, P450, clk ,rst);
VNU_2 VNU451(Q139_451, Q163_451, R139_451, R163_451, L451, P451, clk ,rst);
VNU_2 VNU452(Q140_452, Q164_452, R140_452, R164_452, L452, P452, clk ,rst);
VNU_2 VNU453(Q141_453, Q165_453, R141_453, R165_453, L453, P453, clk ,rst);
VNU_2 VNU454(Q142_454, Q166_454, R142_454, R166_454, L454, P454, clk ,rst);
VNU_2 VNU455(Q143_455, Q167_455, R143_455, R167_455, L455, P455, clk ,rst);
VNU_2 VNU456(Q144_456, Q168_456, R144_456, R168_456, L456, P456, clk ,rst);
VNU_2 VNU457(Q145_457, Q169_457, R145_457, R169_457, L457, P457, clk ,rst);
VNU_2 VNU458(Q146_458, Q170_458, R146_458, R170_458, L458, P458, clk ,rst);
VNU_2 VNU459(Q147_459, Q171_459, R147_459, R171_459, L459, P459, clk ,rst);
VNU_2 VNU460(Q148_460, Q172_460, R148_460, R172_460, L460, P460, clk ,rst);
VNU_2 VNU461(Q149_461, Q173_461, R149_461, R173_461, L461, P461, clk ,rst);
VNU_2 VNU462(Q150_462, Q174_462, R150_462, R174_462, L462, P462, clk ,rst);
VNU_2 VNU463(Q151_463, Q175_463, R151_463, R175_463, L463, P463, clk ,rst);
VNU_2 VNU464(Q152_464, Q176_464, R152_464, R176_464, L464, P464, clk ,rst);
VNU_2 VNU465(Q153_465, Q177_465, R153_465, R177_465, L465, P465, clk ,rst);
VNU_2 VNU466(Q154_466, Q178_466, R154_466, R178_466, L466, P466, clk ,rst);
VNU_2 VNU467(Q155_467, Q179_467, R155_467, R179_467, L467, P467, clk ,rst);
VNU_2 VNU468(Q156_468, Q180_468, R156_468, R180_468, L468, P468, clk ,rst);
VNU_2 VNU469(Q157_469, Q181_469, R157_469, R181_469, L469, P469, clk ,rst);
VNU_2 VNU470(Q158_470, Q182_470, R158_470, R182_470, L470, P470, clk ,rst);
VNU_2 VNU471(Q159_471, Q183_471, R159_471, R183_471, L471, P471, clk ,rst);
VNU_2 VNU472(Q160_472, Q184_472, R160_472, R184_472, L472, P472, clk ,rst);
VNU_2 VNU473(Q161_473, Q185_473, R161_473, R185_473, L473, P473, clk ,rst);
VNU_2 VNU474(Q162_474, Q186_474, R162_474, R186_474, L474, P474, clk ,rst);
VNU_2 VNU475(Q163_475, Q187_475, R163_475, R187_475, L475, P475, clk ,rst);
VNU_2 VNU476(Q164_476, Q188_476, R164_476, R188_476, L476, P476, clk ,rst);
VNU_2 VNU477(Q165_477, Q189_477, R165_477, R189_477, L477, P477, clk ,rst);
VNU_2 VNU478(Q166_478, Q190_478, R166_478, R190_478, L478, P478, clk ,rst);
VNU_2 VNU479(Q167_479, Q191_479, R167_479, R191_479, L479, P479, clk ,rst);
VNU_2 VNU480(Q168_480, Q192_480, R168_480, R192_480, L480, P480, clk ,rst);
VNU_2 VNU481(Q169_481, Q193_481, R169_481, R193_481, L481, P481, clk ,rst);
VNU_2 VNU482(Q170_482, Q194_482, R170_482, R194_482, L482, P482, clk ,rst);
VNU_2 VNU483(Q171_483, Q195_483, R171_483, R195_483, L483, P483, clk ,rst);
VNU_2 VNU484(Q172_484, Q196_484, R172_484, R196_484, L484, P484, clk ,rst);
VNU_2 VNU485(Q173_485, Q197_485, R173_485, R197_485, L485, P485, clk ,rst);
VNU_2 VNU486(Q174_486, Q198_486, R174_486, R198_486, L486, P486, clk ,rst);
VNU_2 VNU487(Q175_487, Q199_487, R175_487, R199_487, L487, P487, clk ,rst);
VNU_2 VNU488(Q176_488, Q200_488, R176_488, R200_488, L488, P488, clk ,rst);
VNU_2 VNU489(Q177_489, Q201_489, R177_489, R201_489, L489, P489, clk ,rst);
VNU_2 VNU490(Q178_490, Q202_490, R178_490, R202_490, L490, P490, clk ,rst);
VNU_2 VNU491(Q179_491, Q203_491, R179_491, R203_491, L491, P491, clk ,rst);
VNU_2 VNU492(Q180_492, Q204_492, R180_492, R204_492, L492, P492, clk ,rst);
VNU_2 VNU493(Q181_493, Q205_493, R181_493, R205_493, L493, P493, clk ,rst);
VNU_2 VNU494(Q182_494, Q206_494, R182_494, R206_494, L494, P494, clk ,rst);
VNU_2 VNU495(Q183_495, Q207_495, R183_495, R207_495, L495, P495, clk ,rst);
VNU_2 VNU496(Q184_496, Q208_496, R184_496, R208_496, L496, P496, clk ,rst);
VNU_2 VNU497(Q185_497, Q209_497, R185_497, R209_497, L497, P497, clk ,rst);
VNU_2 VNU498(Q186_498, Q210_498, R186_498, R210_498, L498, P498, clk ,rst);
VNU_2 VNU499(Q187_499, Q211_499, R187_499, R211_499, L499, P499, clk ,rst);
VNU_2 VNU500(Q188_500, Q212_500, R188_500, R212_500, L500, P500, clk ,rst);
VNU_2 VNU501(Q189_501, Q213_501, R189_501, R213_501, L501, P501, clk ,rst);
VNU_2 VNU502(Q190_502, Q214_502, R190_502, R214_502, L502, P502, clk ,rst);
VNU_2 VNU503(Q191_503, Q215_503, R191_503, R215_503, L503, P503, clk ,rst);
VNU_2 VNU504(Q192_504, Q216_504, R192_504, R216_504, L504, P504, clk ,rst);
VNU_2 VNU505(Q193_505, Q217_505, R193_505, R217_505, L505, P505, clk ,rst);
VNU_2 VNU506(Q194_506, Q218_506, R194_506, R218_506, L506, P506, clk ,rst);
VNU_2 VNU507(Q195_507, Q219_507, R195_507, R219_507, L507, P507, clk ,rst);
VNU_2 VNU508(Q196_508, Q220_508, R196_508, R220_508, L508, P508, clk ,rst);
VNU_2 VNU509(Q197_509, Q221_509, R197_509, R221_509, L509, P509, clk ,rst);
VNU_2 VNU510(Q198_510, Q222_510, R198_510, R222_510, L510, P510, clk ,rst);
VNU_2 VNU511(Q199_511, Q223_511, R199_511, R223_511, L511, P511, clk ,rst);
VNU_2 VNU512(Q200_512, Q224_512, R200_512, R224_512, L512, P512, clk ,rst);
VNU_2 VNU513(Q201_513, Q225_513, R201_513, R225_513, L513, P513, clk ,rst);
VNU_2 VNU514(Q202_514, Q226_514, R202_514, R226_514, L514, P514, clk ,rst);
VNU_2 VNU515(Q203_515, Q227_515, R203_515, R227_515, L515, P515, clk ,rst);
VNU_2 VNU516(Q204_516, Q228_516, R204_516, R228_516, L516, P516, clk ,rst);
VNU_2 VNU517(Q205_517, Q229_517, R205_517, R229_517, L517, P517, clk ,rst);
VNU_2 VNU518(Q206_518, Q230_518, R206_518, R230_518, L518, P518, clk ,rst);
VNU_2 VNU519(Q207_519, Q231_519, R207_519, R231_519, L519, P519, clk ,rst);
VNU_2 VNU520(Q208_520, Q232_520, R208_520, R232_520, L520, P520, clk ,rst);
VNU_2 VNU521(Q209_521, Q233_521, R209_521, R233_521, L521, P521, clk ,rst);
VNU_2 VNU522(Q210_522, Q234_522, R210_522, R234_522, L522, P522, clk ,rst);
VNU_2 VNU523(Q211_523, Q235_523, R211_523, R235_523, L523, P523, clk ,rst);
VNU_2 VNU524(Q212_524, Q236_524, R212_524, R236_524, L524, P524, clk ,rst);
VNU_2 VNU525(Q213_525, Q237_525, R213_525, R237_525, L525, P525, clk ,rst);
VNU_2 VNU526(Q214_526, Q238_526, R214_526, R238_526, L526, P526, clk ,rst);
VNU_2 VNU527(Q215_527, Q239_527, R215_527, R239_527, L527, P527, clk ,rst);
VNU_2 VNU528(Q216_528, Q240_528, R216_528, R240_528, L528, P528, clk ,rst);
VNU_2 VNU529(Q217_529, Q241_529, R217_529, R241_529, L529, P529, clk ,rst);
VNU_2 VNU530(Q218_530, Q242_530, R218_530, R242_530, L530, P530, clk ,rst);
VNU_2 VNU531(Q219_531, Q243_531, R219_531, R243_531, L531, P531, clk ,rst);
VNU_2 VNU532(Q220_532, Q244_532, R220_532, R244_532, L532, P532, clk ,rst);
VNU_2 VNU533(Q221_533, Q245_533, R221_533, R245_533, L533, P533, clk ,rst);
VNU_2 VNU534(Q222_534, Q246_534, R222_534, R246_534, L534, P534, clk ,rst);
VNU_2 VNU535(Q223_535, Q247_535, R223_535, R247_535, L535, P535, clk ,rst);
VNU_2 VNU536(Q224_536, Q248_536, R224_536, R248_536, L536, P536, clk ,rst);
VNU_2 VNU537(Q225_537, Q249_537, R225_537, R249_537, L537, P537, clk ,rst);
VNU_2 VNU538(Q226_538, Q250_538, R226_538, R250_538, L538, P538, clk ,rst);
VNU_2 VNU539(Q227_539, Q251_539, R227_539, R251_539, L539, P539, clk ,rst);
VNU_2 VNU540(Q228_540, Q252_540, R228_540, R252_540, L540, P540, clk ,rst);
VNU_2 VNU541(Q229_541, Q253_541, R229_541, R253_541, L541, P541, clk ,rst);
VNU_2 VNU542(Q230_542, Q254_542, R230_542, R254_542, L542, P542, clk ,rst);
VNU_2 VNU543(Q231_543, Q255_543, R231_543, R255_543, L543, P543, clk ,rst);
VNU_2 VNU544(Q232_544, Q256_544, R232_544, R256_544, L544, P544, clk ,rst);
VNU_2 VNU545(Q233_545, Q257_545, R233_545, R257_545, L545, P545, clk ,rst);
VNU_2 VNU546(Q234_546, Q258_546, R234_546, R258_546, L546, P546, clk ,rst);
VNU_2 VNU547(Q235_547, Q259_547, R235_547, R259_547, L547, P547, clk ,rst);
VNU_2 VNU548(Q236_548, Q260_548, R236_548, R260_548, L548, P548, clk ,rst);
VNU_2 VNU549(Q237_549, Q261_549, R237_549, R261_549, L549, P549, clk ,rst);
VNU_2 VNU550(Q238_550, Q262_550, R238_550, R262_550, L550, P550, clk ,rst);
VNU_2 VNU551(Q239_551, Q263_551, R239_551, R263_551, L551, P551, clk ,rst);
VNU_2 VNU552(Q240_552, Q264_552, R240_552, R264_552, L552, P552, clk ,rst);
VNU_2 VNU553(Q241_553, Q265_553, R241_553, R265_553, L553, P553, clk ,rst);
VNU_2 VNU554(Q242_554, Q266_554, R242_554, R266_554, L554, P554, clk ,rst);
VNU_2 VNU555(Q243_555, Q267_555, R243_555, R267_555, L555, P555, clk ,rst);
VNU_2 VNU556(Q244_556, Q268_556, R244_556, R268_556, L556, P556, clk ,rst);
VNU_2 VNU557(Q245_557, Q269_557, R245_557, R269_557, L557, P557, clk ,rst);
VNU_2 VNU558(Q246_558, Q270_558, R246_558, R270_558, L558, P558, clk ,rst);
VNU_2 VNU559(Q247_559, Q271_559, R247_559, R271_559, L559, P559, clk ,rst);
VNU_2 VNU560(Q248_560, Q272_560, R248_560, R272_560, L560, P560, clk ,rst);
VNU_2 VNU561(Q249_561, Q273_561, R249_561, R273_561, L561, P561, clk ,rst);
VNU_2 VNU562(Q250_562, Q274_562, R250_562, R274_562, L562, P562, clk ,rst);
VNU_2 VNU563(Q251_563, Q275_563, R251_563, R275_563, L563, P563, clk ,rst);
VNU_2 VNU564(Q252_564, Q276_564, R252_564, R276_564, L564, P564, clk ,rst);
VNU_2 VNU565(Q253_565, Q277_565, R253_565, R277_565, L565, P565, clk ,rst);
VNU_2 VNU566(Q254_566, Q278_566, R254_566, R278_566, L566, P566, clk ,rst);
VNU_2 VNU567(Q255_567, Q279_567, R255_567, R279_567, L567, P567, clk ,rst);
VNU_2 VNU568(Q256_568, Q280_568, R256_568, R280_568, L568, P568, clk ,rst);
VNU_2 VNU569(Q257_569, Q281_569, R257_569, R281_569, L569, P569, clk ,rst);
VNU_2 VNU570(Q258_570, Q282_570, R258_570, R282_570, L570, P570, clk ,rst);
VNU_2 VNU571(Q259_571, Q283_571, R259_571, R283_571, L571, P571, clk ,rst);
VNU_2 VNU572(Q260_572, Q284_572, R260_572, R284_572, L572, P572, clk ,rst);
VNU_2 VNU573(Q261_573, Q285_573, R261_573, R285_573, L573, P573, clk ,rst);
VNU_2 VNU574(Q262_574, Q286_574, R262_574, R286_574, L574, P574, clk ,rst);
VNU_2 VNU575(Q263_575, Q287_575, R263_575, R287_575, L575, P575, clk ,rst);
VNU_2 VNU576(Q264_576, Q288_576, R264_576, R288_576, L576, P576, clk ,rst);
endmodule

module VNU_2(
output reg signed [31:0] Q1,
output reg signed [31:0] Q2,
input  signed [31:0] R1,
input  signed [31:0] R2,
input  signed [31:0] L,
output P,
input clk,
input rst);

reg signed [31:0] P_sample;



assign P = P_sample[31] ? 1'b1 : 1'b0;


always@(posedge clk or posedge rst)
begin
if (rst)
begin
Q1 = L;
Q2 = L;
end
else
begin
P_sample = R1 + R2 + L;
Q1 = P_sample - R1;
Q2 = P_sample - R2;
end
end
endmodule

module VNU_3(
output reg signed [31:0] Q1,
output reg signed [31:0] Q2,
output reg signed [31:0] Q3,
input  signed [31:0] R1,
input  signed [31:0] R2,
input  signed [31:0] R3,
input  signed [31:0] L,
output P,
input clk,
input rst);

reg signed [31:0] P_sample;


assign P = P_sample[31] ? 1'b1 : 1'b0;

always@(posedge clk or posedge rst)
begin
if (rst)
begin
Q1 = L;
Q2 = L;
Q3 = L;
end
else
begin
P_sample = R1 + R2 + R3 + L;
Q1 = P_sample - R1;
Q2 = P_sample - R2;
Q3 = P_sample - R3;
end
end

endmodule

module VNU_6(
output reg signed [31:0] Q1,
output reg signed [31:0] Q2,
output reg signed [31:0] Q3,
output reg signed [31:0] Q4,
output reg signed [31:0] Q5,
output reg signed [31:0] Q6,
input  signed [31:0] R1,
input  signed [31:0] R2,
input  signed [31:0] R3,
input  signed [31:0] R4,
input  signed [31:0] R5,
input  signed [31:0] R6,
input  signed [31:0] L,
output P,
input clk,
input rst);

reg signed [31:0] P_sample;



assign P = P_sample[31]? 1'b1 : 1'b0;

always@(posedge clk or posedge rst)
begin

if(rst)
begin
P_sample = L;
Q1 = L;
Q2 = L;
Q3 = L;
Q4 = L;
Q5 = L;
Q6 = L;
end
else
begin
P_sample = R1 + R2 + R3 + R4 + R5 + R6 + L;
Q1 = P_sample - R1;
Q2 = P_sample - R2;
Q3 = P_sample - R3;
Q4 = P_sample - R4;
Q5 = P_sample - R5;
Q6 = P_sample - R6;
end
end
endmodule

module CNU_6(
output reg signed [31:0] R1,
output reg signed [31:0] R2,
output reg signed [31:0] R3,
output reg signed [31:0] R4,
output reg signed [31:0] R5,
output reg signed [31:0] R6,
input signed [31:0] Q1,
input signed [31:0] Q2,
input signed [31:0] Q3,
input signed [31:0] Q4,
input signed [31:0] Q5,
input signed [31:0] Q6,
input clk);

reg signed [31:0] min_sum_1;
reg signed [31:0] min_sum_2;
reg signed [31:0] min_sum_3;
reg signed [31:0] min_sum_4;
reg signed [31:0] min_sum_5;
reg signed [31:0] min_sum_6;
wire [5:0] Q_signs;
wire final_sign_1;
wire final_sign_2;
wire final_sign_3;
wire final_sign_4;
wire final_sign_5;
wire final_sign_6;
wire [31:0] Q1_abs;
wire [31:0] Q2_abs;
wire [31:0] Q3_abs;
wire [31:0] Q4_abs;
wire [31:0] Q5_abs;
wire [31:0] Q6_abs;

assign Q1_abs = (Q1[31]==1) ? ~Q1+1'b1 : Q1;
assign Q2_abs = (Q2[31]==1) ? ~Q2+1'b1 : Q2;
assign Q3_abs = (Q3[31]==1) ? ~Q3+1'b1 : Q3;
assign Q4_abs = (Q4[31]==1) ? ~Q4+1'b1 : Q4;
assign Q5_abs = (Q5[31]==1) ? ~Q5+1'b1 : Q5;
assign Q6_abs = (Q6[31]==1) ? ~Q6+1'b1 : Q6;


assign Q_signs[0] = (Q1[31]==1) ? 1'b1 : 1'b0;
assign Q_signs[1] = (Q2[31]==1) ? 1'b1 : 1'b0;
assign Q_signs[2] = (Q3[31]==1) ? 1'b1 : 1'b0;
assign Q_signs[3] = (Q4[31]==1) ? 1'b1 : 1'b0;
assign Q_signs[4] = (Q5[31]==1) ? 1'b1 : 1'b0;
assign Q_signs[5] = (Q6[31]==1) ? 1'b1 : 1'b0;

assign final_sign_1 = Q_signs[1]^Q_signs[2]^Q_signs[3]^Q_signs[4]^Q_signs[5];
assign final_sign_2 = Q_signs[0]^Q_signs[2]^Q_signs[3]^Q_signs[4]^Q_signs[5];
assign final_sign_3 = Q_signs[1]^Q_signs[0]^Q_signs[3]^Q_signs[4]^Q_signs[5];
assign final_sign_4 = Q_signs[1]^Q_signs[2]^Q_signs[0]^Q_signs[4]^Q_signs[5];
assign final_sign_5 = Q_signs[1]^Q_signs[2]^Q_signs[3]^Q_signs[0]^Q_signs[5];
assign final_sign_6 = Q_signs[1]^Q_signs[2]^Q_signs[3]^Q_signs[4]^Q_signs[0];



always@(negedge clk)
begin

if (Q2_abs<=Q3_abs && Q2_abs<=Q4_abs && Q2_abs<=Q5_abs && Q2_abs<=Q6_abs) begin min_sum_1 = Q2_abs;  end 
if (Q3_abs<Q2_abs  && Q3_abs<=Q4_abs && Q3_abs<=Q5_abs && Q3_abs<=Q6_abs) begin min_sum_1 = Q3_abs;  end 
if (Q4_abs<Q2_abs  && Q4_abs<Q3_abs && Q4_abs<=Q5_abs && Q4_abs<=Q6_abs)  begin min_sum_1 = Q4_abs;  end
if (Q5_abs<Q2_abs  && Q5_abs<Q3_abs && Q5_abs<Q4_abs && Q5_abs<=Q6_abs)   begin min_sum_1 = Q5_abs;  end 
if (Q6_abs<Q2_abs  && Q6_abs<Q3_abs && Q6_abs<Q4_abs && Q6_abs<Q5_abs )   begin min_sum_1 = Q6_abs;  end 

if (Q1_abs<=Q3_abs && Q1_abs<=Q4_abs && Q1_abs<=Q5_abs && Q1_abs<=Q6_abs) begin min_sum_2 = Q1_abs;  end 
if (Q3_abs<Q1_abs  && Q3_abs<=Q4_abs && Q3_abs<=Q5_abs && Q3_abs<=Q6_abs) begin min_sum_2 = Q3_abs;  end 
if (Q4_abs<Q1_abs  && Q4_abs<Q3_abs && Q4_abs<=Q5_abs && Q4_abs<=Q6_abs)  begin min_sum_2 = Q4_abs;  end
if (Q5_abs<Q1_abs  && Q5_abs<Q3_abs && Q5_abs<Q4_abs && Q5_abs<=Q6_abs)   begin min_sum_2 = Q5_abs;  end 
if (Q6_abs<Q1_abs  && Q6_abs<Q3_abs && Q6_abs<Q4_abs && Q6_abs<Q5_abs )   begin min_sum_2 = Q6_abs;  end 

if (Q2_abs<=Q1_abs && Q2_abs<=Q4_abs && Q2_abs<=Q5_abs && Q2_abs<=Q6_abs) begin min_sum_3 = Q2_abs;  end 
if (Q1_abs<Q2_abs  && Q1_abs<=Q4_abs && Q1_abs<=Q5_abs && Q1_abs<=Q6_abs) begin min_sum_3 = Q1_abs;  end 
if (Q4_abs<Q2_abs  && Q4_abs<Q1_abs && Q4_abs<=Q5_abs && Q4_abs<=Q6_abs)  begin min_sum_3 = Q4_abs;  end
if (Q5_abs<Q2_abs  && Q5_abs<Q1_abs && Q5_abs<Q4_abs && Q5_abs<=Q6_abs)   begin min_sum_3 = Q5_abs;  end 
if (Q6_abs<Q2_abs  && Q6_abs<Q1_abs && Q6_abs<Q4_abs && Q6_abs<Q5_abs )   begin min_sum_3 = Q6_abs;  end 

if (Q2_abs<=Q3_abs && Q2_abs<=Q1_abs && Q2_abs<=Q5_abs && Q2_abs<=Q6_abs) begin min_sum_4 = Q2_abs;  end 
if (Q3_abs<Q2_abs  && Q3_abs<=Q1_abs && Q3_abs<=Q5_abs && Q3_abs<=Q6_abs) begin min_sum_4 = Q3_abs;  end 
if (Q1_abs<Q2_abs  && Q1_abs<Q3_abs && Q1_abs<=Q5_abs && Q1_abs<=Q6_abs)  begin min_sum_4 = Q1_abs;  end
if (Q5_abs<Q2_abs  && Q5_abs<Q3_abs && Q5_abs<Q1_abs && Q5_abs<=Q6_abs)   begin min_sum_4 = Q5_abs;  end 
if (Q6_abs<Q2_abs  && Q6_abs<Q3_abs && Q6_abs<Q1_abs && Q6_abs<Q5_abs )   begin min_sum_4 = Q6_abs;  end 

if (Q2_abs<=Q3_abs && Q2_abs<=Q4_abs && Q2_abs<=Q1_abs && Q2_abs<=Q6_abs) begin min_sum_5 = Q2_abs;  end 
if (Q3_abs<Q2_abs  && Q3_abs<=Q4_abs && Q3_abs<=Q1_abs && Q3_abs<=Q6_abs) begin min_sum_5 = Q3_abs;  end 
if (Q4_abs<Q2_abs  && Q4_abs<Q3_abs && Q4_abs<=Q1_abs && Q4_abs<=Q6_abs)  begin min_sum_5 = Q4_abs;  end
if (Q1_abs<Q2_abs  && Q1_abs<Q3_abs && Q1_abs<Q4_abs && Q1_abs<=Q6_abs)   begin min_sum_5 = Q1_abs;  end 
if (Q6_abs<Q2_abs  && Q6_abs<Q3_abs && Q6_abs<Q4_abs && Q6_abs<Q1_abs )   begin min_sum_5 = Q6_abs;  end 

if (Q2_abs<=Q3_abs && Q2_abs<=Q4_abs && Q2_abs<=Q5_abs && Q2_abs<=Q1_abs) begin min_sum_6 = Q2_abs;  end 
if (Q3_abs<Q2_abs  && Q3_abs<=Q4_abs && Q3_abs<=Q5_abs && Q3_abs<=Q1_abs) begin min_sum_6 = Q3_abs;  end 
if (Q4_abs<Q2_abs  && Q4_abs<Q3_abs && Q4_abs<=Q5_abs && Q4_abs<=Q1_abs)  begin min_sum_6 = Q4_abs;  end
if (Q5_abs<Q2_abs  && Q5_abs<Q3_abs && Q5_abs<Q4_abs && Q5_abs<=Q1_abs)   begin min_sum_6 = Q5_abs;  end 
if (Q1_abs<Q2_abs  && Q1_abs<Q3_abs && Q1_abs<Q4_abs && Q1_abs<Q5_abs )   begin min_sum_6 = Q1_abs;  end 

R1 = final_sign_1 ? ~min_sum_1 + 1'b1 : min_sum_1;
R2 = final_sign_2 ? ~min_sum_2 + 1'b1 : min_sum_2;
R3 = final_sign_3 ? ~min_sum_3 + 1'b1 : min_sum_3;
R4 = final_sign_4 ? ~min_sum_4 + 1'b1 : min_sum_4;
R5 = final_sign_5 ? ~min_sum_5 + 1'b1 : min_sum_5;
R6 = final_sign_6 ? ~min_sum_6 + 1'b1 : min_sum_6;

end

endmodule

module CNU_7(
output reg signed [31:0] R1,
output reg signed [31:0] R2,
output reg signed [31:0] R3,
output reg signed [31:0] R4,
output reg signed [31:0] R5,
output reg signed [31:0] R6,
output reg signed [31:0] R7,
input signed [31:0] Q1,
input signed [31:0] Q2,
input signed [31:0] Q3,
input signed [31:0] Q4,
input signed [31:0] Q5,
input signed [31:0] Q6,
input signed [31:0] Q7,
input clk);

reg signed [31:0] min_sum_1;
reg signed [31:0] min_sum_2;
reg signed [31:0] min_sum_3;
reg signed [31:0] min_sum_4;
reg signed [31:0] min_sum_5;
reg signed [31:0] min_sum_6;
reg signed [31:0] min_sum_7;
wire [6:0] Q_signs;
wire final_sign_1;
wire final_sign_2;
wire final_sign_3;
wire final_sign_4;
wire final_sign_5;
wire final_sign_6;
wire final_sign_7;
wire [31:0] Q1_abs;
wire [31:0] Q2_abs;
wire [31:0] Q3_abs;
wire [31:0] Q4_abs;
wire [31:0] Q5_abs;
wire [31:0] Q6_abs;
wire [31:0] Q7_abs;

assign Q1_abs = (Q1[31]==1) ? ~Q1+1'b1 : Q1;
assign Q2_abs = (Q2[31]==1) ? ~Q2+1'b1 : Q2;
assign Q3_abs = (Q3[31]==1) ? ~Q3+1'b1 : Q3;
assign Q4_abs = (Q4[31]==1) ? ~Q4+1'b1 : Q4;
assign Q5_abs = (Q5[31]==1) ? ~Q5+1'b1 : Q5;
assign Q6_abs = (Q6[31]==1) ? ~Q6+1'b1 : Q6;
assign Q7_abs = (Q7[31]==1) ? ~Q7+1'b1 : Q7;


assign Q_signs[0] = (Q1[31]==1) ? 1'b1 : 1'b0;
assign Q_signs[1] = (Q2[31]==1) ? 1'b1 : 1'b0;
assign Q_signs[2] = (Q3[31]==1) ? 1'b1 : 1'b0;
assign Q_signs[3] = (Q4[31]==1) ? 1'b1 : 1'b0;
assign Q_signs[4] = (Q5[31]==1) ? 1'b1 : 1'b0;
assign Q_signs[5] = (Q6[31]==1) ? 1'b1 : 1'b0;
assign Q_signs[6] = (Q7[31]==1) ? 1'b1 : 1'b0;

assign final_sign_1 = Q_signs[1]^Q_signs[2]^Q_signs[3]^Q_signs[4]^Q_signs[5]^Q_signs[6];
assign final_sign_2 = Q_signs[0]^Q_signs[2]^Q_signs[3]^Q_signs[4]^Q_signs[5]^Q_signs[6];
assign final_sign_3 = Q_signs[1]^Q_signs[0]^Q_signs[3]^Q_signs[4]^Q_signs[5]^Q_signs[6];
assign final_sign_4 = Q_signs[1]^Q_signs[2]^Q_signs[0]^Q_signs[4]^Q_signs[5]^Q_signs[6];
assign final_sign_5 = Q_signs[1]^Q_signs[2]^Q_signs[3]^Q_signs[0]^Q_signs[5]^Q_signs[6];
assign final_sign_6 = Q_signs[1]^Q_signs[2]^Q_signs[3]^Q_signs[4]^Q_signs[0]^Q_signs[6];
assign final_sign_7 = Q_signs[1]^Q_signs[2]^Q_signs[3]^Q_signs[4]^Q_signs[5]^Q_signs[0];


always@(negedge clk)
begin

if (Q2_abs<=Q3_abs && Q2_abs<=Q4_abs && Q2_abs<=Q5_abs && Q2_abs<=Q6_abs && Q2_abs<=Q7_abs) begin min_sum_1 = Q2_abs;  end 
if (Q3_abs<Q2_abs  && Q3_abs<=Q4_abs && Q3_abs<=Q5_abs && Q3_abs<=Q6_abs && Q3_abs<=Q7_abs) begin min_sum_1 = Q3_abs;  end 
if (Q4_abs<Q2_abs  && Q4_abs<Q3_abs && Q4_abs<=Q5_abs && Q4_abs<=Q6_abs && Q4_abs<=Q7_abs)  begin min_sum_1 = Q4_abs;  end
if (Q5_abs<Q2_abs  && Q5_abs<Q3_abs && Q5_abs<Q4_abs && Q5_abs<=Q6_abs && Q5_abs<=Q7_abs)   begin min_sum_1 = Q5_abs;  end 
if (Q6_abs<Q2_abs  && Q6_abs<Q3_abs && Q6_abs<Q4_abs && Q6_abs<Q5_abs  && Q6_abs<=Q7_abs)   begin min_sum_1 = Q6_abs;  end 
if (Q7_abs<Q2_abs  && Q7_abs<Q3_abs && Q7_abs<Q4_abs && Q7_abs<Q5_abs  && Q7_abs<=Q6_abs)   begin min_sum_1 = Q7_abs;  end 

if (Q1_abs<=Q3_abs && Q1_abs<=Q4_abs && Q1_abs<=Q5_abs && Q1_abs<=Q6_abs && Q1_abs<=Q7_abs) begin min_sum_2 = Q1_abs;  end 
if (Q3_abs<Q1_abs  && Q3_abs<=Q4_abs && Q3_abs<=Q5_abs && Q3_abs<=Q6_abs && Q3_abs<=Q7_abs) begin min_sum_2 = Q3_abs;  end 
if (Q4_abs<Q1_abs  && Q4_abs<Q3_abs && Q4_abs<=Q5_abs && Q4_abs<=Q6_abs && Q4_abs<=Q7_abs)  begin min_sum_2 = Q4_abs;  end
if (Q5_abs<Q1_abs  && Q5_abs<Q3_abs && Q5_abs<Q4_abs && Q5_abs<=Q6_abs && Q5_abs<=Q7_abs)   begin min_sum_2 = Q5_abs;  end 
if (Q6_abs<Q1_abs  && Q6_abs<Q3_abs && Q6_abs<Q4_abs && Q6_abs<Q5_abs  && Q6_abs<=Q7_abs)   begin min_sum_2 = Q6_abs;  end 
if (Q7_abs<Q1_abs  && Q7_abs<Q3_abs && Q7_abs<Q4_abs && Q7_abs<Q5_abs  && Q7_abs<=Q6_abs)   begin min_sum_2 = Q7_abs;  end 

if (Q2_abs<=Q1_abs && Q2_abs<=Q4_abs && Q2_abs<=Q5_abs && Q2_abs<=Q6_abs && Q2_abs<=Q7_abs) begin min_sum_3 = Q2_abs;  end 
if (Q1_abs<Q2_abs  && Q1_abs<=Q4_abs && Q1_abs<=Q5_abs && Q1_abs<=Q6_abs && Q1_abs<=Q7_abs) begin min_sum_3 = Q1_abs;  end 
if (Q4_abs<Q2_abs  && Q4_abs<Q1_abs && Q4_abs<=Q5_abs && Q4_abs<=Q6_abs && Q4_abs<=Q7_abs)  begin min_sum_3 = Q4_abs;  end
if (Q5_abs<Q2_abs  && Q5_abs<Q1_abs && Q5_abs<Q4_abs && Q5_abs<=Q6_abs && Q5_abs<=Q7_abs)   begin min_sum_3 = Q5_abs;  end 
if (Q6_abs<Q2_abs  && Q6_abs<Q1_abs && Q6_abs<Q4_abs && Q6_abs<Q5_abs  && Q6_abs<=Q7_abs)   begin min_sum_3 = Q6_abs;  end 
if (Q7_abs<Q2_abs  && Q7_abs<Q1_abs && Q7_abs<Q4_abs && Q7_abs<Q5_abs  && Q7_abs<=Q6_abs)   begin min_sum_3 = Q7_abs;  end 

if (Q2_abs<=Q3_abs && Q2_abs<=Q1_abs && Q2_abs<=Q5_abs && Q2_abs<=Q6_abs && Q2_abs<=Q7_abs) begin min_sum_4 = Q2_abs;  end 
if (Q3_abs<Q2_abs  && Q3_abs<=Q1_abs && Q3_abs<=Q5_abs && Q3_abs<=Q6_abs && Q3_abs<=Q7_abs) begin min_sum_4 = Q3_abs;  end 
if (Q1_abs<Q2_abs  && Q1_abs<Q3_abs && Q1_abs<=Q5_abs && Q1_abs<=Q6_abs && Q1_abs<=Q7_abs)  begin min_sum_4 = Q1_abs;  end
if (Q5_abs<Q2_abs  && Q5_abs<Q3_abs && Q5_abs<Q1_abs && Q5_abs<=Q6_abs && Q5_abs<=Q7_abs)   begin min_sum_4 = Q5_abs;  end 
if (Q6_abs<Q2_abs  && Q6_abs<Q3_abs && Q6_abs<Q1_abs && Q6_abs<Q5_abs && Q6_abs<=Q7_abs )   begin min_sum_4 = Q6_abs;  end 
if (Q7_abs<Q2_abs  && Q7_abs<Q3_abs && Q7_abs<Q1_abs && Q7_abs<Q5_abs  && Q7_abs<=Q6_abs)   begin min_sum_4 = Q7_abs;  end 

if (Q2_abs<=Q3_abs && Q2_abs<=Q4_abs && Q2_abs<=Q1_abs && Q2_abs<=Q6_abs && Q2_abs<=Q7_abs) begin min_sum_5 = Q2_abs;  end 
if (Q3_abs<Q2_abs  && Q3_abs<=Q4_abs && Q3_abs<=Q1_abs && Q3_abs<=Q6_abs && Q3_abs<=Q7_abs) begin min_sum_5 = Q3_abs;  end 
if (Q4_abs<Q2_abs  && Q4_abs<Q3_abs && Q4_abs<=Q1_abs && Q4_abs<=Q6_abs && Q4_abs<=Q7_abs)  begin min_sum_5 = Q4_abs;  end
if (Q1_abs<Q2_abs  && Q1_abs<Q3_abs && Q1_abs<Q4_abs && Q1_abs<=Q6_abs && Q1_abs<=Q7_abs)   begin min_sum_5 = Q1_abs;  end 
if (Q6_abs<Q2_abs  && Q6_abs<Q3_abs && Q6_abs<Q4_abs && Q6_abs<Q1_abs  && Q6_abs<=Q7_abs)   begin min_sum_5 = Q6_abs;  end 
if (Q7_abs<Q2_abs  && Q7_abs<Q3_abs && Q7_abs<Q4_abs && Q7_abs<Q1_abs  && Q7_abs<=Q6_abs)   begin min_sum_5 = Q7_abs;  end 

if (Q2_abs<=Q3_abs && Q2_abs<=Q4_abs && Q2_abs<=Q5_abs && Q2_abs<=Q1_abs && Q2_abs<=Q7_abs) begin min_sum_6 = Q2_abs;  end 
if (Q3_abs<Q2_abs  && Q3_abs<=Q4_abs && Q3_abs<=Q5_abs && Q3_abs<=Q1_abs && Q3_abs<=Q7_abs) begin min_sum_6 = Q3_abs;  end 
if (Q4_abs<Q2_abs  && Q4_abs<Q3_abs && Q4_abs<=Q5_abs && Q4_abs<=Q1_abs && Q4_abs<=Q7_abs)  begin min_sum_6 = Q4_abs;  end
if (Q5_abs<Q2_abs  && Q5_abs<Q3_abs && Q5_abs<Q4_abs && Q5_abs<=Q1_abs && Q5_abs<=Q7_abs)   begin min_sum_6 = Q5_abs;  end 
if (Q1_abs<Q2_abs  && Q1_abs<Q3_abs && Q1_abs<Q4_abs && Q1_abs<Q5_abs  && Q1_abs<=Q7_abs)   begin min_sum_6 = Q1_abs;  end 
if (Q7_abs<Q2_abs  && Q7_abs<Q3_abs && Q7_abs<Q4_abs && Q7_abs<Q5_abs  && Q7_abs<=Q1_abs)   begin min_sum_6 = Q7_abs;  end 

if (Q2_abs<=Q3_abs && Q2_abs<=Q4_abs && Q2_abs<=Q5_abs && Q2_abs<=Q1_abs && Q2_abs<=Q6_abs) begin min_sum_7 = Q2_abs;  end 
if (Q3_abs<Q2_abs  && Q3_abs<=Q4_abs && Q3_abs<=Q5_abs && Q3_abs<=Q1_abs && Q3_abs<=Q6_abs) begin min_sum_7 = Q3_abs;  end 
if (Q4_abs<Q2_abs  && Q4_abs<Q3_abs && Q4_abs<=Q5_abs && Q4_abs<=Q1_abs && Q4_abs<=Q6_abs)  begin min_sum_7 = Q4_abs;  end
if (Q5_abs<Q2_abs  && Q5_abs<Q3_abs && Q5_abs<Q4_abs && Q5_abs<=Q1_abs && Q5_abs<=Q6_abs)   begin min_sum_7 = Q5_abs;  end 
if (Q1_abs<Q2_abs  && Q1_abs<Q3_abs && Q1_abs<Q4_abs && Q1_abs<Q5_abs  && Q1_abs<=Q6_abs)   begin min_sum_7 = Q1_abs;  end 
if (Q6_abs<Q2_abs  && Q6_abs<Q3_abs && Q6_abs<Q4_abs && Q6_abs<Q5_abs  && Q6_abs<=Q1_abs)   begin min_sum_7 = Q6_abs;  end 

R1 = final_sign_1 ? ~min_sum_1 + 1'b1 : min_sum_1;
R2 = final_sign_2 ? ~min_sum_2 + 1'b1 : min_sum_2;
R3 = final_sign_3 ? ~min_sum_3 + 1'b1 : min_sum_3;
R4 = final_sign_4 ? ~min_sum_4 + 1'b1 : min_sum_4;
R5 = final_sign_5 ? ~min_sum_5 + 1'b1 : min_sum_5;
R6 = final_sign_6 ? ~min_sum_6 + 1'b1 : min_sum_6;
R7 = final_sign_7 ? ~min_sum_7 + 1'b1 : min_sum_7;

end

endmodule